`timescale 1us / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:57:26 11/16/2015 
// Design Name: 
// Module Name:    fir400 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 401 tap FIR filter
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fir400( // 27 MHz clock, ready asserted with frequency of 48 kHz
  input wire clock,reset,ready,
  input wire signed [9:0] coeff,
  input wire signed [17:0] x,
  output wire signed [17:0] y,
  output reg [8:0] index
);

	reg signed [17:0] audio_out;
	assign y = audio_out;
	reg signed [27:0] accumulator; 
	reg signed [17:0] sample [511:0];  // 512 element array each 8 bits wide
	reg [8:0] offset = 0; // increment offset with each sample to always point to the newest sample
	
	always @(posedge clock) begin
		if (reset == 1) begin
			accumulator <= 0;
			index <= 0;
			offset <= 0;
		end
		else if (ready == 1) begin // reset accumulator to begin calculations for new audio sample
			accumulator <= 0;
			offset <= offset +1; 
			index <= 0;
			sample[(offset+1) & 5'b1111_1] <= x;
		end
// 		pipeline to perform FIR 401-tap filter multiplication and addition over 401 cycles 
		else if (index<401) begin 
			accumulator <= accumulator + coeff*sample[(offset-index)& 5'b1111_1]; // delay 1
			index <= index + 1;
		end
		else begin
			audio_out <= accumulator[27:10];
		end
		
	end
endmodule

//////////////////////////////////////////////////////////////////////////////////////////
/// coefficients for the 401-tap FIR filters stored in ROM for the various filters
//////////////////////////////////////////////////////////////////////////////////////////


module coeffs400tap_test(
  input wire [8:0] index,
  output reg signed [9:0] coeff
);
  // tools will turn this into a 400x10 ROM
  always @(index)
    case (index)
		9'd0:  coeff = 10'sd0; 
		9'd1:  coeff = 10'sd0; 
		9'd2:  coeff = 10'sd0; 
		9'd3:  coeff = 10'sd0; 
		9'd4:  coeff = 10'sd0; 
		9'd5:  coeff = 10'sd0; 
		9'd6:  coeff = 10'sd0; 
		9'd7:  coeff = 10'sd0; 
		9'd8:  coeff = 10'sd0; 
		9'd9:  coeff = 10'sd0; 
		9'd10:  coeff = 10'sd0; 
		9'd11:  coeff = 10'sd0; 
		9'd12:  coeff = 10'sd0; 
		9'd13:  coeff = 10'sd0; 
		9'd14:  coeff = 10'sd0; 
		9'd15:  coeff = 10'sd0; 
		9'd16:  coeff = 10'sd0; 
		9'd17:  coeff = 10'sd0; 
		9'd18:  coeff = 10'sd0; 
		9'd19:  coeff = 10'sd0; 
		9'd20:  coeff = 10'sd0; 
		9'd21:  coeff = 10'sd0; 
		9'd22:  coeff = 10'sd0; 
		9'd23:  coeff = 10'sd0; 
		9'd24:  coeff = 10'sd0; 
		9'd25:  coeff = 10'sd0; 
		9'd26:  coeff = 10'sd0; 
		9'd27:  coeff = 10'sd0; 
		9'd28:  coeff = 10'sd0; 
		9'd29:  coeff = 10'sd0; 
		9'd30:  coeff = 10'sd0; 
		9'd31:  coeff = 10'sd0; 
		9'd32:  coeff = 10'sd0; 
		9'd33:  coeff = 10'sd0; 
		9'd34:  coeff = 10'sd0; 
		9'd35:  coeff = 10'sd0; 
		9'd36:  coeff = 10'sd0; 
		9'd37:  coeff = 10'sd0; 
		9'd38:  coeff = 10'sd0; 
		9'd39:  coeff = 10'sd0; 
		9'd40:  coeff = 10'sd0; 
		9'd41:  coeff = 10'sd0; 
		9'd42:  coeff = 10'sd0; 
		9'd43:  coeff = 10'sd0; 
		9'd44:  coeff = 10'sd0; 
		9'd45:  coeff = 10'sd0; 
		9'd46:  coeff = 10'sd0; 
		9'd47:  coeff = 10'sd0; 
		9'd48:  coeff = 10'sd0; 
		9'd49:  coeff = 10'sd0; 
		9'd50:  coeff = 10'sd0; 
		9'd51:  coeff = 10'sd0; 
		9'd52:  coeff = 10'sd0; 
		9'd53:  coeff = 10'sd0; 
		9'd54:  coeff = 10'sd0; 
		9'd55:  coeff = 10'sd0; 
		9'd56:  coeff = 10'sd0; 
		9'd57:  coeff = 10'sd0; 
		9'd58:  coeff = 10'sd0; 
		9'd59:  coeff = 10'sd0; 
		9'd60:  coeff = 10'sd0; 
		9'd61:  coeff = 10'sd0; 
		9'd62:  coeff = 10'sd0; 
		9'd63:  coeff = 10'sd0; 
		9'd64:  coeff = 10'sd0; 
		9'd65:  coeff = 10'sd0; 
		9'd66:  coeff = 10'sd0; 
		9'd67:  coeff = 10'sd0; 
		9'd68:  coeff = 10'sd0; 
		9'd69:  coeff = 10'sd0; 
		9'd70:  coeff = 10'sd0; 
		9'd71:  coeff = 10'sd0; 
		9'd72:  coeff = 10'sd0; 
		9'd73:  coeff = 10'sd0; 
		9'd74:  coeff = 10'sd0; 
		9'd75:  coeff = 10'sd0; 
		9'd76:  coeff = 10'sd0; 
		9'd77:  coeff = 10'sd0; 
		9'd78:  coeff = 10'sd0; 
		9'd79:  coeff = 10'sd0; 
		9'd80:  coeff = 10'sd0; 
		9'd81:  coeff = 10'sd0; 
		9'd82:  coeff = 10'sd0; 
		9'd83:  coeff = 10'sd0; 
		9'd84:  coeff = 10'sd0; 
		9'd85:  coeff = 10'sd0; 
		9'd86:  coeff = 10'sd0; 
		9'd87:  coeff = 10'sd0; 
		9'd88:  coeff = 10'sd0; 
		9'd89:  coeff = 10'sd0; 
		9'd90:  coeff = 10'sd0; 
		9'd91:  coeff = 10'sd0; 
		9'd92:  coeff = 10'sd0; 
		9'd93:  coeff = 10'sd0; 
		9'd94:  coeff = 10'sd0; 
		9'd95:  coeff = 10'sd0; 
		9'd96:  coeff = 10'sd0; 
		9'd97:  coeff = 10'sd0; 
		9'd98:  coeff = 10'sd0; 
		9'd99:  coeff = 10'sd0; 
		9'd100:  coeff = 10'sd0; 
		9'd101:  coeff = 10'sd0; 
		9'd102:  coeff = 10'sd0; 
		9'd103:  coeff = 10'sd0; 
		9'd104:  coeff = 10'sd0; 
		9'd105:  coeff = 10'sd0; 
		9'd106:  coeff = 10'sd0; 
		9'd107:  coeff = 10'sd0; 
		9'd108:  coeff = 10'sd0; 
		9'd109:  coeff = 10'sd0; 
		9'd110:  coeff = 10'sd0; 
		9'd111:  coeff = 10'sd0; 
		9'd112:  coeff = 10'sd0; 
		9'd113:  coeff = 10'sd0; 
		9'd114:  coeff = 10'sd0; 
		9'd115:  coeff = 10'sd0; 
		9'd116:  coeff = 10'sd0; 
		9'd117:  coeff = 10'sd0; 
		9'd118:  coeff = 10'sd0; 
		9'd119:  coeff = 10'sd0; 
		9'd120:  coeff = 10'sd0; 
		9'd121:  coeff = 10'sd0; 
		9'd122:  coeff = 10'sd0; 
		9'd123:  coeff = 10'sd0; 
		9'd124:  coeff = 10'sd0; 
		9'd125:  coeff = 10'sd0; 
		9'd126:  coeff = 10'sd0; 
		9'd127:  coeff = 10'sd0; 
		9'd128:  coeff = 10'sd0; 
		9'd129:  coeff = 10'sd0; 
		9'd130:  coeff = 10'sd0; 
		9'd131:  coeff = 10'sd0; 
		9'd132:  coeff = 10'sd0; 
		9'd133:  coeff = 10'sd0; 
		9'd134:  coeff = 10'sd0; 
		9'd135:  coeff = 10'sd0; 
		9'd136:  coeff = 10'sd0; 
		9'd137:  coeff = 10'sd0; 
		9'd138:  coeff = 10'sd0; 
		9'd139:  coeff = 10'sd0; 
		9'd140:  coeff = 10'sd0; 
		9'd141:  coeff = 10'sd0; 
		9'd142:  coeff = 10'sd0; 
		9'd143:  coeff = 10'sd0; 
		9'd144:  coeff = 10'sd0; 
		9'd145:  coeff = 10'sd0; 
		9'd146:  coeff = 10'sd0; 
		9'd147:  coeff = 10'sd0; 
		9'd148:  coeff = 10'sd0; 
		9'd149:  coeff = 10'sd0; 
		9'd150:  coeff = 10'sd0; 
		9'd151:  coeff = 10'sd0; 
		9'd152:  coeff = 10'sd0; 
		9'd153:  coeff = 10'sd0; 
		9'd154:  coeff = 10'sd0; 
		9'd155:  coeff = 10'sd0; 
		9'd156:  coeff = 10'sd0; 
		9'd157:  coeff = 10'sd0; 
		9'd158:  coeff = 10'sd0; 
		9'd159:  coeff = 10'sd0; 
		9'd160:  coeff = 10'sd0; 
		9'd161:  coeff = 10'sd0; 
		9'd162:  coeff = 10'sd0; 
		9'd163:  coeff = 10'sd0; 
		9'd164:  coeff = 10'sd0; 
		9'd165:  coeff = 10'sd0; 
		9'd166:  coeff = 10'sd0; 
		9'd167:  coeff = 10'sd0; 
		9'd168:  coeff = 10'sd0; 
		9'd169:  coeff = 10'sd0; 
		9'd170:  coeff = 10'sd0; 
		9'd171:  coeff = 10'sd0; 
		9'd172:  coeff = 10'sd0; 
		9'd173:  coeff = 10'sd0; 
		9'd174:  coeff = 10'sd0; 
		9'd175:  coeff = 10'sd0; 
		9'd176:  coeff = 10'sd0; 
		9'd177:  coeff = 10'sd0; 
		9'd178:  coeff = 10'sd0; 
		9'd179:  coeff = 10'sd0; 
		9'd180:  coeff = 10'sd0; 
		9'd181:  coeff = 10'sd0; 
		9'd182:  coeff = 10'sd0; 
		9'd183:  coeff = 10'sd0; 
		9'd184:  coeff = 10'sd0; 
		9'd185:  coeff = 10'sd0; 
		9'd186:  coeff = 10'sd0; 
		9'd187:  coeff = 10'sd0; 
		9'd188:  coeff = 10'sd0; 
		9'd189:  coeff = 10'sd0; 
		9'd190:  coeff = 10'sd0; 
		9'd191:  coeff = 10'sd0; 
		9'd192:  coeff = 10'sd0; 
		9'd193:  coeff = 10'sd0; 
		9'd194:  coeff = 10'sd0; 
		9'd195:  coeff = 10'sd0; 
		9'd196:  coeff = 10'sd0; 
		9'd197:  coeff = 10'sd0; 
		9'd198:  coeff = 10'sd0; 
		9'd199:  coeff = 10'sd0; 
		9'd200:  coeff = 10'sd0; 
		9'd201:  coeff = 10'sd0; 
		9'd202:  coeff = 10'sd0; 
		9'd203:  coeff = 10'sd0; 
		9'd204:  coeff = 10'sd0; 
		9'd205:  coeff = 10'sd0; 
		9'd206:  coeff = 10'sd0; 
		9'd207:  coeff = 10'sd0; 
		9'd208:  coeff = 10'sd0; 
		9'd209:  coeff = 10'sd0; 
		9'd210:  coeff = 10'sd0; 
		9'd211:  coeff = 10'sd0; 
		9'd212:  coeff = 10'sd0; 
		9'd213:  coeff = 10'sd0; 
		9'd214:  coeff = 10'sd0; 
		9'd215:  coeff = 10'sd0; 
		9'd216:  coeff = 10'sd0; 
		9'd217:  coeff = 10'sd0; 
		9'd218:  coeff = 10'sd0; 
		9'd219:  coeff = 10'sd0; 
		9'd220:  coeff = 10'sd0; 
		9'd221:  coeff = 10'sd0; 
		9'd222:  coeff = 10'sd0; 
		9'd223:  coeff = 10'sd0; 
		9'd224:  coeff = 10'sd0; 
		9'd225:  coeff = 10'sd0; 
		9'd226:  coeff = 10'sd0; 
		9'd227:  coeff = 10'sd0; 
		9'd228:  coeff = 10'sd0; 
		9'd229:  coeff = 10'sd0; 
		9'd230:  coeff = 10'sd0; 
		9'd231:  coeff = 10'sd0; 
		9'd232:  coeff = 10'sd0; 
		9'd233:  coeff = 10'sd0; 
		9'd234:  coeff = 10'sd0; 
		9'd235:  coeff = 10'sd0; 
		9'd236:  coeff = 10'sd0; 
		9'd237:  coeff = 10'sd0; 
		9'd238:  coeff = 10'sd0; 
		9'd239:  coeff = 10'sd0; 
		9'd240:  coeff = 10'sd0; 
		9'd241:  coeff = 10'sd0; 
		9'd242:  coeff = 10'sd0; 
		9'd243:  coeff = 10'sd0; 
		9'd244:  coeff = 10'sd0; 
		9'd245:  coeff = 10'sd0; 
		9'd246:  coeff = 10'sd0; 
		9'd247:  coeff = 10'sd0; 
		9'd248:  coeff = 10'sd0; 
		9'd249:  coeff = 10'sd0; 
		9'd250:  coeff = 10'sd0; 
		9'd251:  coeff = 10'sd0; 
		9'd252:  coeff = 10'sd0; 
		9'd253:  coeff = 10'sd0; 
		9'd254:  coeff = 10'sd0; 
		9'd255:  coeff = 10'sd0; 
		9'd256:  coeff = 10'sd0; 
		9'd257:  coeff = 10'sd0; 
		9'd258:  coeff = 10'sd0; 
		9'd259:  coeff = 10'sd0; 
		9'd260:  coeff = 10'sd0; 
		9'd261:  coeff = 10'sd0; 
		9'd262:  coeff = 10'sd0; 
		9'd263:  coeff = 10'sd0; 
		9'd264:  coeff = 10'sd0; 
		9'd265:  coeff = 10'sd0; 
		9'd266:  coeff = 10'sd0; 
		9'd267:  coeff = 10'sd0; 
		9'd268:  coeff = 10'sd0; 
		9'd269:  coeff = 10'sd0; 
		9'd270:  coeff = 10'sd0; 
		9'd271:  coeff = 10'sd0; 
		9'd272:  coeff = 10'sd0; 
		9'd273:  coeff = 10'sd0; 
		9'd274:  coeff = 10'sd0; 
		9'd275:  coeff = 10'sd0; 
		9'd276:  coeff = 10'sd0; 
		9'd277:  coeff = 10'sd0; 
		9'd278:  coeff = 10'sd0; 
		9'd279:  coeff = 10'sd0; 
		9'd280:  coeff = 10'sd0; 
		9'd281:  coeff = 10'sd0; 
		9'd282:  coeff = 10'sd0; 
		9'd283:  coeff = 10'sd0; 
		9'd284:  coeff = 10'sd0; 
		9'd285:  coeff = 10'sd0; 
		9'd286:  coeff = 10'sd0; 
		9'd287:  coeff = 10'sd0; 
		9'd288:  coeff = 10'sd0; 
		9'd289:  coeff = 10'sd0; 
		9'd290:  coeff = 10'sd0; 
		9'd291:  coeff = 10'sd0; 
		9'd292:  coeff = 10'sd0; 
		9'd293:  coeff = 10'sd0; 
		9'd294:  coeff = 10'sd0; 
		9'd295:  coeff = 10'sd0; 
		9'd296:  coeff = 10'sd0; 
		9'd297:  coeff = 10'sd0; 
		9'd298:  coeff = 10'sd0; 
		9'd299:  coeff = 10'sd0; 
		9'd300:  coeff = 10'sd0; 
		9'd301:  coeff = 10'sd0; 
		9'd302:  coeff = 10'sd0; 
		9'd303:  coeff = 10'sd0; 
		9'd304:  coeff = 10'sd0; 
		9'd305:  coeff = 10'sd0; 
		9'd306:  coeff = 10'sd0; 
		9'd307:  coeff = 10'sd0; 
		9'd308:  coeff = 10'sd0; 
		9'd309:  coeff = 10'sd0; 
		9'd310:  coeff = 10'sd0; 
		9'd311:  coeff = 10'sd0; 
		9'd312:  coeff = 10'sd0; 
		9'd313:  coeff = 10'sd0; 
		9'd314:  coeff = 10'sd0; 
		9'd315:  coeff = 10'sd0; 
		9'd316:  coeff = 10'sd0; 
		9'd317:  coeff = 10'sd0; 
		9'd318:  coeff = 10'sd0; 
		9'd319:  coeff = 10'sd0; 
		9'd320:  coeff = 10'sd0; 
		9'd321:  coeff = 10'sd0; 
		9'd322:  coeff = 10'sd0; 
		9'd323:  coeff = 10'sd0; 
		9'd324:  coeff = 10'sd0; 
		9'd325:  coeff = 10'sd0; 
		9'd326:  coeff = 10'sd0; 
		9'd327:  coeff = 10'sd0; 
		9'd328:  coeff = 10'sd0; 
		9'd329:  coeff = 10'sd0; 
		9'd330:  coeff = 10'sd0; 
		9'd331:  coeff = 10'sd0; 
		9'd332:  coeff = 10'sd0; 
		9'd333:  coeff = 10'sd0; 
		9'd334:  coeff = 10'sd0; 
		9'd335:  coeff = 10'sd0; 
		9'd336:  coeff = 10'sd0; 
		9'd337:  coeff = 10'sd0; 
		9'd338:  coeff = 10'sd0; 
		9'd339:  coeff = 10'sd0; 
		9'd340:  coeff = 10'sd0; 
		9'd341:  coeff = 10'sd0; 
		9'd342:  coeff = 10'sd0; 
		9'd343:  coeff = 10'sd0; 
		9'd344:  coeff = 10'sd0; 
		9'd345:  coeff = 10'sd0; 
		9'd346:  coeff = 10'sd0; 
		9'd347:  coeff = 10'sd0; 
		9'd348:  coeff = 10'sd0; 
		9'd349:  coeff = 10'sd0; 
		9'd350:  coeff = 10'sd0; 
		9'd351:  coeff = 10'sd0; 
		9'd352:  coeff = 10'sd0; 
		9'd353:  coeff = 10'sd0; 
		9'd354:  coeff = 10'sd0; 
		9'd355:  coeff = 10'sd0; 
		9'd356:  coeff = 10'sd0; 
		9'd357:  coeff = 10'sd0; 
		9'd358:  coeff = 10'sd0; 
		9'd359:  coeff = 10'sd0; 
		9'd360:  coeff = 10'sd0; 
		9'd361:  coeff = 10'sd0; 
		9'd362:  coeff = 10'sd0; 
		9'd363:  coeff = 10'sd0; 
		9'd364:  coeff = 10'sd0; 
		9'd365:  coeff = 10'sd0; 
		9'd366:  coeff = 10'sd0; 
		9'd367:  coeff = 10'sd0; 
		9'd368:  coeff = 10'sd0; 
		9'd369:  coeff = 10'sd0; 
		9'd370:  coeff = 10'sd0; 
		9'd371:  coeff = 10'sd0; 
		9'd372:  coeff = 10'sd0; 
		9'd373:  coeff = 10'sd0; 
		9'd374:  coeff = 10'sd0; 
		9'd375:  coeff = 10'sd0; 
		9'd376:  coeff = 10'sd0; 
		9'd377:  coeff = 10'sd0; 
		9'd378:  coeff = 10'sd0; 
		9'd379:  coeff = 10'sd0; 
		9'd380:  coeff = 10'sd0; 
		9'd381:  coeff = 10'sd0; 
		9'd382:  coeff = 10'sd0; 
		9'd383:  coeff = 10'sd0; 
		9'd384:  coeff = 10'sd0; 
		9'd385:  coeff = 10'sd0; 
		9'd386:  coeff = 10'sd0; 
		9'd387:  coeff = 10'sd0; 
		9'd388:  coeff = 10'sd0; 
		9'd389:  coeff = 10'sd0; 
		9'd390:  coeff = 10'sd0; 
		9'd391:  coeff = 10'sd0; 
		9'd392:  coeff = 10'sd0; 
		9'd393:  coeff = 10'sd0; 
		9'd394:  coeff = 10'sd0; 
		9'd395:  coeff = 10'sd0; 
		9'd396:  coeff = 10'sd0; 
		9'd397:  coeff = 10'sd0; 
		9'd398:  coeff = 10'sd0; 
		9'd399:  coeff = 10'sd0; 
		9'd400:  coeff = 10'sd511; 
	 
      default: coeff = 10'hXXX;
    endcase
endmodule

	 

module coeffs400tap_below120Hz(
  input wire [8:0] index,
  output reg signed [9:0] coeff
);
  // tools will turn this into a 400x10 ROM
  always @(index)
    case (index)

		9'd0:  coeff = 10'sd0; 
		9'd1:  coeff = 10'sd0; 
		9'd2:  coeff = 10'sd0; 
		9'd3:  coeff = 10'sd0; 
		9'd4:  coeff = 10'sd0; 
		9'd5:  coeff = 10'sd0; 
		9'd6:  coeff = 10'sd0; 
		9'd7:  coeff = 10'sd0; 
		9'd8:  coeff = 10'sd0; 
		9'd9:  coeff = 10'sd0; 
		9'd10:  coeff = 10'sd0; 
		9'd11:  coeff = 10'sd0; 
		9'd12:  coeff = 10'sd0; 
		9'd13:  coeff = 10'sd0; 
		9'd14:  coeff = 10'sd0; 
		9'd15:  coeff = 10'sd0; 
		9'd16:  coeff = 10'sd0; 
		9'd17:  coeff = 10'sd0; 
		9'd18:  coeff = 10'sd0; 
		9'd19:  coeff = 10'sd0; 
		9'd20:  coeff = 10'sd0; 
		9'd21:  coeff = 10'sd0; 
		9'd22:  coeff = 10'sd0; 
		9'd23:  coeff = 10'sd0; 
		9'd24:  coeff = 10'sd0; 
		9'd25:  coeff = 10'sd0; 
		9'd26:  coeff = 10'sd0; 
		9'd27:  coeff = 10'sd0; 
		9'd28:  coeff = 10'sd0; 
		9'd29:  coeff = 10'sd0; 
		9'd30:  coeff = 10'sd0; 
		9'd31:  coeff = 10'sd0; 
		9'd32:  coeff = 10'sd0; 
		9'd33:  coeff = 10'sd0; 
		9'd34:  coeff = 10'sd0; 
		9'd35:  coeff = 10'sd0; 
		9'd36:  coeff = 10'sd0; 
		9'd37:  coeff = 10'sd0; 
		9'd38:  coeff = 10'sd0; 
		9'd39:  coeff = 10'sd0; 
		9'd40:  coeff = 10'sd0; 
		9'd41:  coeff = 10'sd0; 
		9'd42:  coeff = 10'sd0; 
		9'd43:  coeff = 10'sd0; 
		9'd44:  coeff = 10'sd0; 
		9'd45:  coeff = 10'sd0; 
		9'd46:  coeff = 10'sd0; 
		9'd47:  coeff = 10'sd0; 
		9'd48:  coeff = 10'sd0; 
		9'd49:  coeff = 10'sd0; 
		9'd50:  coeff = 10'sd0; 
		9'd51:  coeff = 10'sd0; 
		9'd52:  coeff = 10'sd0; 
		9'd53:  coeff = 10'sd0; 
		9'd54:  coeff = 10'sd0; 
		9'd55:  coeff = 10'sd0; 
		9'd56:  coeff = 10'sd0; 
		9'd57:  coeff = 10'sd0; 
		9'd58:  coeff = 10'sd0; 
		9'd59:  coeff = 10'sd0; 
		9'd60:  coeff = 10'sd0; 
		9'd61:  coeff = 10'sd0; 
		9'd62:  coeff = 10'sd0; 
		9'd63:  coeff = 10'sd0; 
		9'd64:  coeff = 10'sd0; 
		9'd65:  coeff = 10'sd0; 
		9'd66:  coeff = 10'sd0; 
		9'd67:  coeff = 10'sd0; 
		9'd68:  coeff = 10'sd0; 
		9'd69:  coeff = 10'sd0; 
		9'd70:  coeff = 10'sd0; 
		9'd71:  coeff = 10'sd0; 
		9'd72:  coeff = 10'sd0; 
		9'd73:  coeff = 10'sd0; 
		9'd74:  coeff = 10'sd0; 
		9'd75:  coeff = 10'sd0; 
		9'd76:  coeff = 10'sd0; 
		9'd77:  coeff = 10'sd0; 
		9'd78:  coeff = 10'sd0; 
		9'd79:  coeff = 10'sd0; 
		9'd80:  coeff = 10'sd0; 
		9'd81:  coeff = 10'sd1; 
		9'd82:  coeff = 10'sd1; 
		9'd83:  coeff = 10'sd1; 
		9'd84:  coeff = 10'sd1; 
		9'd85:  coeff = 10'sd1; 
		9'd86:  coeff = 10'sd1; 
		9'd87:  coeff = 10'sd1; 
		9'd88:  coeff = 10'sd1; 
		9'd89:  coeff = 10'sd1; 
		9'd90:  coeff = 10'sd1; 
		9'd91:  coeff = 10'sd1; 
		9'd92:  coeff = 10'sd1; 
		9'd93:  coeff = 10'sd1; 
		9'd94:  coeff = 10'sd1; 
		9'd95:  coeff = 10'sd1; 
		9'd96:  coeff = 10'sd1; 
		9'd97:  coeff = 10'sd1; 
		9'd98:  coeff = 10'sd1; 
		9'd99:  coeff = 10'sd1; 
		9'd100:  coeff = 10'sd1; 
		9'd101:  coeff = 10'sd1; 
		9'd102:  coeff = 10'sd1; 
		9'd103:  coeff = 10'sd1; 
		9'd104:  coeff = 10'sd1; 
		9'd105:  coeff = 10'sd1; 
		9'd106:  coeff = 10'sd2; 
		9'd107:  coeff = 10'sd2; 
		9'd108:  coeff = 10'sd2; 
		9'd109:  coeff = 10'sd2; 
		9'd110:  coeff = 10'sd2; 
		9'd111:  coeff = 10'sd2; 
		9'd112:  coeff = 10'sd2; 
		9'd113:  coeff = 10'sd2; 
		9'd114:  coeff = 10'sd2; 
		9'd115:  coeff = 10'sd2; 
		9'd116:  coeff = 10'sd2; 
		9'd117:  coeff = 10'sd2; 
		9'd118:  coeff = 10'sd2; 
		9'd119:  coeff = 10'sd2; 
		9'd120:  coeff = 10'sd2; 
		9'd121:  coeff = 10'sd3; 
		9'd122:  coeff = 10'sd3; 
		9'd123:  coeff = 10'sd3; 
		9'd124:  coeff = 10'sd3; 
		9'd125:  coeff = 10'sd3; 
		9'd126:  coeff = 10'sd3; 
		9'd127:  coeff = 10'sd3; 
		9'd128:  coeff = 10'sd3; 
		9'd129:  coeff = 10'sd3; 
		9'd130:  coeff = 10'sd3; 
		9'd131:  coeff = 10'sd3; 
		9'd132:  coeff = 10'sd3; 
		9'd133:  coeff = 10'sd3; 
		9'd134:  coeff = 10'sd4; 
		9'd135:  coeff = 10'sd4; 
		9'd136:  coeff = 10'sd4; 
		9'd137:  coeff = 10'sd4; 
		9'd138:  coeff = 10'sd4; 
		9'd139:  coeff = 10'sd4; 
		9'd140:  coeff = 10'sd4; 
		9'd141:  coeff = 10'sd4; 
		9'd142:  coeff = 10'sd4; 
		9'd143:  coeff = 10'sd4; 
		9'd144:  coeff = 10'sd4; 
		9'd145:  coeff = 10'sd5; 
		9'd146:  coeff = 10'sd5; 
		9'd147:  coeff = 10'sd5; 
		9'd148:  coeff = 10'sd5; 
		9'd149:  coeff = 10'sd5; 
		9'd150:  coeff = 10'sd5; 
		9'd151:  coeff = 10'sd5; 
		9'd152:  coeff = 10'sd5; 
		9'd153:  coeff = 10'sd5; 
		9'd154:  coeff = 10'sd5; 
		9'd155:  coeff = 10'sd5; 
		9'd156:  coeff = 10'sd6; 
		9'd157:  coeff = 10'sd6; 
		9'd158:  coeff = 10'sd6; 
		9'd159:  coeff = 10'sd6; 
		9'd160:  coeff = 10'sd6; 
		9'd161:  coeff = 10'sd6; 
		9'd162:  coeff = 10'sd6; 
		9'd163:  coeff = 10'sd6; 
		9'd164:  coeff = 10'sd6; 
		9'd165:  coeff = 10'sd6; 
		9'd166:  coeff = 10'sd6; 
		9'd167:  coeff = 10'sd6; 
		9'd168:  coeff = 10'sd7; 
		9'd169:  coeff = 10'sd7; 
		9'd170:  coeff = 10'sd7; 
		9'd171:  coeff = 10'sd7; 
		9'd172:  coeff = 10'sd7; 
		9'd173:  coeff = 10'sd7; 
		9'd174:  coeff = 10'sd7; 
		9'd175:  coeff = 10'sd7; 
		9'd176:  coeff = 10'sd7; 
		9'd177:  coeff = 10'sd7; 
		9'd178:  coeff = 10'sd7; 
		9'd179:  coeff = 10'sd7; 
		9'd180:  coeff = 10'sd7; 
		9'd181:  coeff = 10'sd7; 
		9'd182:  coeff = 10'sd7; 
		9'd183:  coeff = 10'sd7; 
		9'd184:  coeff = 10'sd8; 
		9'd185:  coeff = 10'sd8; 
		9'd186:  coeff = 10'sd8; 
		9'd187:  coeff = 10'sd8; 
		9'd188:  coeff = 10'sd8; 
		9'd189:  coeff = 10'sd8; 
		9'd190:  coeff = 10'sd8; 
		9'd191:  coeff = 10'sd8; 
		9'd192:  coeff = 10'sd8; 
		9'd193:  coeff = 10'sd8; 
		9'd194:  coeff = 10'sd8; 
		9'd195:  coeff = 10'sd8; 
		9'd196:  coeff = 10'sd8; 
		9'd197:  coeff = 10'sd8; 
		9'd198:  coeff = 10'sd8; 
		9'd199:  coeff = 10'sd8; 
		9'd200:  coeff = 10'sd8; 
		9'd201:  coeff = 10'sd8; 
		9'd202:  coeff = 10'sd8; 
		9'd203:  coeff = 10'sd8; 
		9'd204:  coeff = 10'sd8; 
		9'd205:  coeff = 10'sd8; 
		9'd206:  coeff = 10'sd8; 
		9'd207:  coeff = 10'sd8; 
		9'd208:  coeff = 10'sd8; 
		9'd209:  coeff = 10'sd8; 
		9'd210:  coeff = 10'sd8; 
		9'd211:  coeff = 10'sd8; 
		9'd212:  coeff = 10'sd8; 
		9'd213:  coeff = 10'sd8; 
		9'd214:  coeff = 10'sd8; 
		9'd215:  coeff = 10'sd8; 
		9'd216:  coeff = 10'sd8; 
		9'd217:  coeff = 10'sd7; 
		9'd218:  coeff = 10'sd7; 
		9'd219:  coeff = 10'sd7; 
		9'd220:  coeff = 10'sd7; 
		9'd221:  coeff = 10'sd7; 
		9'd222:  coeff = 10'sd7; 
		9'd223:  coeff = 10'sd7; 
		9'd224:  coeff = 10'sd7; 
		9'd225:  coeff = 10'sd7; 
		9'd226:  coeff = 10'sd7; 
		9'd227:  coeff = 10'sd7; 
		9'd228:  coeff = 10'sd7; 
		9'd229:  coeff = 10'sd7; 
		9'd230:  coeff = 10'sd7; 
		9'd231:  coeff = 10'sd7; 
		9'd232:  coeff = 10'sd7; 
		9'd233:  coeff = 10'sd6; 
		9'd234:  coeff = 10'sd6; 
		9'd235:  coeff = 10'sd6; 
		9'd236:  coeff = 10'sd6; 
		9'd237:  coeff = 10'sd6; 
		9'd238:  coeff = 10'sd6; 
		9'd239:  coeff = 10'sd6; 
		9'd240:  coeff = 10'sd6; 
		9'd241:  coeff = 10'sd6; 
		9'd242:  coeff = 10'sd6; 
		9'd243:  coeff = 10'sd6; 
		9'd244:  coeff = 10'sd6; 
		9'd245:  coeff = 10'sd5; 
		9'd246:  coeff = 10'sd5; 
		9'd247:  coeff = 10'sd5; 
		9'd248:  coeff = 10'sd5; 
		9'd249:  coeff = 10'sd5; 
		9'd250:  coeff = 10'sd5; 
		9'd251:  coeff = 10'sd5; 
		9'd252:  coeff = 10'sd5; 
		9'd253:  coeff = 10'sd5; 
		9'd254:  coeff = 10'sd5; 
		9'd255:  coeff = 10'sd5; 
		9'd256:  coeff = 10'sd4; 
		9'd257:  coeff = 10'sd4; 
		9'd258:  coeff = 10'sd4; 
		9'd259:  coeff = 10'sd4; 
		9'd260:  coeff = 10'sd4; 
		9'd261:  coeff = 10'sd4; 
		9'd262:  coeff = 10'sd4; 
		9'd263:  coeff = 10'sd4; 
		9'd264:  coeff = 10'sd4; 
		9'd265:  coeff = 10'sd4; 
		9'd266:  coeff = 10'sd4; 
		9'd267:  coeff = 10'sd3; 
		9'd268:  coeff = 10'sd3; 
		9'd269:  coeff = 10'sd3; 
		9'd270:  coeff = 10'sd3; 
		9'd271:  coeff = 10'sd3; 
		9'd272:  coeff = 10'sd3; 
		9'd273:  coeff = 10'sd3; 
		9'd274:  coeff = 10'sd3; 
		9'd275:  coeff = 10'sd3; 
		9'd276:  coeff = 10'sd3; 
		9'd277:  coeff = 10'sd3; 
		9'd278:  coeff = 10'sd3; 
		9'd279:  coeff = 10'sd3; 
		9'd280:  coeff = 10'sd2; 
		9'd281:  coeff = 10'sd2; 
		9'd282:  coeff = 10'sd2; 
		9'd283:  coeff = 10'sd2; 
		9'd284:  coeff = 10'sd2; 
		9'd285:  coeff = 10'sd2; 
		9'd286:  coeff = 10'sd2; 
		9'd287:  coeff = 10'sd2; 
		9'd288:  coeff = 10'sd2; 
		9'd289:  coeff = 10'sd2; 
		9'd290:  coeff = 10'sd2; 
		9'd291:  coeff = 10'sd2; 
		9'd292:  coeff = 10'sd2; 
		9'd293:  coeff = 10'sd2; 
		9'd294:  coeff = 10'sd2; 
		9'd295:  coeff = 10'sd1; 
		9'd296:  coeff = 10'sd1; 
		9'd297:  coeff = 10'sd1; 
		9'd298:  coeff = 10'sd1; 
		9'd299:  coeff = 10'sd1; 
		9'd300:  coeff = 10'sd1; 
		9'd301:  coeff = 10'sd1; 
		9'd302:  coeff = 10'sd1; 
		9'd303:  coeff = 10'sd1; 
		9'd304:  coeff = 10'sd1; 
		9'd305:  coeff = 10'sd1; 
		9'd306:  coeff = 10'sd1; 
		9'd307:  coeff = 10'sd1; 
		9'd308:  coeff = 10'sd1; 
		9'd309:  coeff = 10'sd1; 
		9'd310:  coeff = 10'sd1; 
		9'd311:  coeff = 10'sd1; 
		9'd312:  coeff = 10'sd1; 
		9'd313:  coeff = 10'sd1; 
		9'd314:  coeff = 10'sd1; 
		9'd315:  coeff = 10'sd1; 
		9'd316:  coeff = 10'sd1; 
		9'd317:  coeff = 10'sd1; 
		9'd318:  coeff = 10'sd1; 
		9'd319:  coeff = 10'sd1; 
		9'd320:  coeff = 10'sd0; 
		9'd321:  coeff = 10'sd0; 
		9'd322:  coeff = 10'sd0; 
		9'd323:  coeff = 10'sd0; 
		9'd324:  coeff = 10'sd0; 
		9'd325:  coeff = 10'sd0; 
		9'd326:  coeff = 10'sd0; 
		9'd327:  coeff = 10'sd0; 
		9'd328:  coeff = 10'sd0; 
		9'd329:  coeff = 10'sd0; 
		9'd330:  coeff = 10'sd0; 
		9'd331:  coeff = 10'sd0; 
		9'd332:  coeff = 10'sd0; 
		9'd333:  coeff = 10'sd0; 
		9'd334:  coeff = 10'sd0; 
		9'd335:  coeff = 10'sd0; 
		9'd336:  coeff = 10'sd0; 
		9'd337:  coeff = 10'sd0; 
		9'd338:  coeff = 10'sd0; 
		9'd339:  coeff = 10'sd0; 
		9'd340:  coeff = 10'sd0; 
		9'd341:  coeff = 10'sd0; 
		9'd342:  coeff = 10'sd0; 
		9'd343:  coeff = 10'sd0; 
		9'd344:  coeff = 10'sd0; 
		9'd345:  coeff = 10'sd0; 
		9'd346:  coeff = 10'sd0; 
		9'd347:  coeff = 10'sd0; 
		9'd348:  coeff = 10'sd0; 
		9'd349:  coeff = 10'sd0; 
		9'd350:  coeff = 10'sd0; 
		9'd351:  coeff = 10'sd0; 
		9'd352:  coeff = 10'sd0; 
		9'd353:  coeff = 10'sd0; 
		9'd354:  coeff = 10'sd0; 
		9'd355:  coeff = 10'sd0; 
		9'd356:  coeff = 10'sd0; 
		9'd357:  coeff = 10'sd0; 
		9'd358:  coeff = 10'sd0; 
		9'd359:  coeff = 10'sd0; 
		9'd360:  coeff = 10'sd0; 
		9'd361:  coeff = 10'sd0; 
		9'd362:  coeff = 10'sd0; 
		9'd363:  coeff = 10'sd0; 
		9'd364:  coeff = 10'sd0; 
		9'd365:  coeff = 10'sd0; 
		9'd366:  coeff = 10'sd0; 
		9'd367:  coeff = 10'sd0; 
		9'd368:  coeff = 10'sd0; 
		9'd369:  coeff = 10'sd0; 
		9'd370:  coeff = 10'sd0; 
		9'd371:  coeff = 10'sd0; 
		9'd372:  coeff = 10'sd0; 
		9'd373:  coeff = 10'sd0; 
		9'd374:  coeff = 10'sd0; 
		9'd375:  coeff = 10'sd0; 
		9'd376:  coeff = 10'sd0; 
		9'd377:  coeff = 10'sd0; 
		9'd378:  coeff = 10'sd0; 
		9'd379:  coeff = 10'sd0; 
		9'd380:  coeff = 10'sd0; 
		9'd381:  coeff = 10'sd0; 
		9'd382:  coeff = 10'sd0; 
		9'd383:  coeff = 10'sd0; 
		9'd384:  coeff = 10'sd0; 
		9'd385:  coeff = 10'sd0; 
		9'd386:  coeff = 10'sd0; 
		9'd387:  coeff = 10'sd0; 
		9'd388:  coeff = 10'sd0; 
		9'd389:  coeff = 10'sd0; 
		9'd390:  coeff = 10'sd0; 
		9'd391:  coeff = 10'sd0; 
		9'd392:  coeff = 10'sd0; 
		9'd393:  coeff = 10'sd0; 
		9'd394:  coeff = 10'sd0; 
		9'd395:  coeff = 10'sd0; 
		9'd396:  coeff = 10'sd0; 
		9'd397:  coeff = 10'sd0; 
		9'd398:  coeff = 10'sd0; 
		9'd399:  coeff = 10'sd0; 
		9'd400:  coeff = 10'sd0; 

      default: coeff = 10'hXXX;
    endcase
endmodule

// not the best way to build an all pass filter
module coeffs_allpass(
  input wire [8:0] index,
  output reg signed [9:0] coeff
);
  // tools will turn this into a 400x10 ROM
	always @(index)
		case (index)
	 
	 
			9'd0:  coeff = 10'sd0; 
			9'd1:  coeff = 10'sd0; 
			9'd2:  coeff = 10'sd0; 
			9'd3:  coeff = 10'sd0; 
			9'd4:  coeff = 10'sd0; 
			9'd5:  coeff = 10'sd0; 
			9'd6:  coeff = 10'sd0; 
			9'd7:  coeff = 10'sd0; 
			9'd8:  coeff = 10'sd0; 
			9'd9:  coeff = 10'sd0; 
			9'd10:  coeff = 10'sd0; 
			9'd11:  coeff = 10'sd0; 
			9'd12:  coeff = 10'sd0; 
			9'd13:  coeff = 10'sd0; 
			9'd14:  coeff = 10'sd0; 
			9'd15:  coeff = 10'sd0; 
			9'd16:  coeff = 10'sd0; 
			9'd17:  coeff = 10'sd0; 
			9'd18:  coeff = 10'sd0; 
			9'd19:  coeff = 10'sd0; 
			9'd20:  coeff = 10'sd0; 
			9'd21:  coeff = 10'sd0; 
			9'd22:  coeff = 10'sd0; 
			9'd23:  coeff = 10'sd0; 
			9'd24:  coeff = 10'sd0; 
			9'd25:  coeff = 10'sd0; 
			9'd26:  coeff = 10'sd0; 
			9'd27:  coeff = 10'sd0; 
			9'd28:  coeff = 10'sd0; 
			9'd29:  coeff = 10'sd0; 
			9'd30:  coeff = 10'sd0; 
			9'd31:  coeff = 10'sd0; 
			9'd32:  coeff = 10'sd0; 
			9'd33:  coeff = 10'sd0; 
			9'd34:  coeff = 10'sd0; 
			9'd35:  coeff = 10'sd0; 
			9'd36:  coeff = 10'sd0; 
			9'd37:  coeff = 10'sd0; 
			9'd38:  coeff = 10'sd0; 
			9'd39:  coeff = 10'sd0; 
			9'd40:  coeff = 10'sd0; 
			9'd41:  coeff = 10'sd0; 
			9'd42:  coeff = 10'sd0; 
			9'd43:  coeff = 10'sd0; 
			9'd44:  coeff = 10'sd0; 
			9'd45:  coeff = 10'sd0; 
			9'd46:  coeff = 10'sd0; 
			9'd47:  coeff = 10'sd0; 
			9'd48:  coeff = 10'sd0; 
			9'd49:  coeff = 10'sd0; 
			9'd50:  coeff = 10'sd0; 
			9'd51:  coeff = 10'sd0; 
			9'd52:  coeff = 10'sd0; 
			9'd53:  coeff = 10'sd0; 
			9'd54:  coeff = 10'sd0; 
			9'd55:  coeff = 10'sd0; 
			9'd56:  coeff = 10'sd0; 
			9'd57:  coeff = 10'sd0; 
			9'd58:  coeff = 10'sd0; 
			9'd59:  coeff = 10'sd0; 
			9'd60:  coeff = 10'sd0; 
			9'd61:  coeff = 10'sd0; 
			9'd62:  coeff = 10'sd0; 
			9'd63:  coeff = 10'sd0; 
			9'd64:  coeff = 10'sd0; 
			9'd65:  coeff = 10'sd0; 
			9'd66:  coeff = 10'sd0; 
			9'd67:  coeff = 10'sd0; 
			9'd68:  coeff = 10'sd0; 
			9'd69:  coeff = 10'sd0; 
			9'd70:  coeff = 10'sd0; 
			9'd71:  coeff = 10'sd0; 
			9'd72:  coeff = 10'sd0; 
			9'd73:  coeff = 10'sd0; 
			9'd74:  coeff = 10'sd0; 
			9'd75:  coeff = 10'sd0; 
			9'd76:  coeff = 10'sd0; 
			9'd77:  coeff = 10'sd0; 
			9'd78:  coeff = 10'sd0; 
			9'd79:  coeff = 10'sd0; 
			9'd80:  coeff = 10'sd0; 
			9'd81:  coeff = 10'sd0; 
			9'd82:  coeff = 10'sd0; 
			9'd83:  coeff = 10'sd0; 
			9'd84:  coeff = 10'sd0; 
			9'd85:  coeff = 10'sd0; 
			9'd86:  coeff = 10'sd0; 
			9'd87:  coeff = 10'sd0; 
			9'd88:  coeff = 10'sd0; 
			9'd89:  coeff = 10'sd0; 
			9'd90:  coeff = 10'sd0; 
			9'd91:  coeff = 10'sd0; 
			9'd92:  coeff = 10'sd0; 
			9'd93:  coeff = 10'sd0; 
			9'd94:  coeff = -10'sd1; 
			9'd95:  coeff = 10'sd1; 
			9'd96:  coeff = -10'sd1; 
			9'd97:  coeff = 10'sd1; 
			9'd98:  coeff = 10'sd0; 
			9'd99:  coeff = 10'sd0; 
			9'd100:  coeff = 10'sd0; 
			9'd101:  coeff = 10'sd0; 
			9'd102:  coeff = 10'sd0; 
			9'd103:  coeff = -10'sd1; 
			9'd104:  coeff = 10'sd1; 
			9'd105:  coeff = -10'sd1; 
			9'd106:  coeff = 10'sd1; 
			9'd107:  coeff = -10'sd1; 
			9'd108:  coeff = 10'sd1; 
			9'd109:  coeff = 10'sd0; 
			9'd110:  coeff = 10'sd0; 
			9'd111:  coeff = 10'sd0; 
			9'd112:  coeff = -10'sd1; 
			9'd113:  coeff = 10'sd1; 
			9'd114:  coeff = -10'sd1; 
			9'd115:  coeff = 10'sd1; 
			9'd116:  coeff = -10'sd1; 
			9'd117:  coeff = 10'sd1; 
			9'd118:  coeff = -10'sd1; 
			9'd119:  coeff = 10'sd0; 
			9'd120:  coeff = 10'sd0; 
			9'd121:  coeff = -10'sd1; 
			9'd122:  coeff = 10'sd1; 
			9'd123:  coeff = -10'sd2; 
			9'd124:  coeff = 10'sd2; 
			9'd125:  coeff = -10'sd2; 
			9'd126:  coeff = 10'sd2; 
			9'd127:  coeff = -10'sd2; 
			9'd128:  coeff = 10'sd1; 
			9'd129:  coeff = -10'sd1; 
			9'd130:  coeff = 10'sd0; 
			9'd131:  coeff = 10'sd1; 
			9'd132:  coeff = -10'sd1; 
			9'd133:  coeff = 10'sd2; 
			9'd134:  coeff = -10'sd3; 
			9'd135:  coeff = 10'sd3; 
			9'd136:  coeff = -10'sd3; 
			9'd137:  coeff = 10'sd2; 
			9'd138:  coeff = -10'sd2; 
			9'd139:  coeff = 10'sd1; 
			9'd140:  coeff = 10'sd0; 
			9'd141:  coeff = -10'sd1; 
			9'd142:  coeff = 10'sd2; 
			9'd143:  coeff = -10'sd3; 
			9'd144:  coeff = 10'sd4; 
			9'd145:  coeff = -10'sd4; 
			9'd146:  coeff = 10'sd4; 
			9'd147:  coeff = -10'sd3; 
			9'd148:  coeff = 10'sd3; 
			9'd149:  coeff = -10'sd1; 
			9'd150:  coeff = 10'sd0; 
			9'd151:  coeff = 10'sd1; 
			9'd152:  coeff = -10'sd3; 
			9'd153:  coeff = 10'sd4; 
			9'd154:  coeff = -10'sd5; 
			9'd155:  coeff = 10'sd6; 
			9'd156:  coeff = -10'sd5; 
			9'd157:  coeff = 10'sd5; 
			9'd158:  coeff = -10'sd4; 
			9'd159:  coeff = 10'sd2; 
			9'd160:  coeff = 10'sd0; 
			9'd161:  coeff = -10'sd2; 
			9'd162:  coeff = 10'sd4; 
			9'd163:  coeff = -10'sd6; 
			9'd164:  coeff = 10'sd7; 
			9'd165:  coeff = -10'sd8; 
			9'd166:  coeff = 10'sd8; 
			9'd167:  coeff = -10'sd7; 
			9'd168:  coeff = 10'sd5; 
			9'd169:  coeff = -10'sd3; 
			9'd170:  coeff = 10'sd0; 
			9'd171:  coeff = 10'sd3; 
			9'd172:  coeff = -10'sd6; 
			9'd173:  coeff = 10'sd9; 
			9'd174:  coeff = -10'sd11; 
			9'd175:  coeff = 10'sd12; 
			9'd176:  coeff = -10'sd12; 
			9'd177:  coeff = 10'sd11; 
			9'd178:  coeff = -10'sd8; 
			9'd179:  coeff = 10'sd5; 
			9'd180:  coeff = 10'sd0; 
			9'd181:  coeff = -10'sd5; 
			9'd182:  coeff = 10'sd10; 
			9'd183:  coeff = -10'sd15; 
			9'd184:  coeff = 10'sd19; 
			9'd185:  coeff = -10'sd21; 
			9'd186:  coeff = 10'sd22; 
			9'd187:  coeff = -10'sd20; 
			9'd188:  coeff = 10'sd16; 
			9'd189:  coeff = -10'sd9; 
			9'd190:  coeff = 10'sd0; 
			9'd191:  coeff = 10'sd11; 
			9'd192:  coeff = -10'sd24; 
			9'd193:  coeff = 10'sd37; 
			9'd194:  coeff = -10'sd51; 
			9'd195:  coeff = 10'sd65; 
			9'd196:  coeff = -10'sd77; 
			9'd197:  coeff = 10'sd88; 
			9'd198:  coeff = -10'sd96; 
			9'd199:  coeff = 10'sd101; 
			9'd200:  coeff = 10'sd922; 
			9'd201:  coeff = 10'sd101; 
			9'd202:  coeff = -10'sd96; 
			9'd203:  coeff = 10'sd88; 
			9'd204:  coeff = -10'sd77; 
			9'd205:  coeff = 10'sd65; 
			9'd206:  coeff = -10'sd51; 
			9'd207:  coeff = 10'sd37; 
			9'd208:  coeff = -10'sd24; 
			9'd209:  coeff = 10'sd11; 
			9'd210:  coeff = 10'sd0; 
			9'd211:  coeff = -10'sd9; 
			9'd212:  coeff = 10'sd16; 
			9'd213:  coeff = -10'sd20; 
			9'd214:  coeff = 10'sd22; 
			9'd215:  coeff = -10'sd21; 
			9'd216:  coeff = 10'sd19; 
			9'd217:  coeff = -10'sd15; 
			9'd218:  coeff = 10'sd10; 
			9'd219:  coeff = -10'sd5; 
			9'd220:  coeff = 10'sd0; 
			9'd221:  coeff = 10'sd5; 
			9'd222:  coeff = -10'sd8; 
			9'd223:  coeff = 10'sd11; 
			9'd224:  coeff = -10'sd12; 
			9'd225:  coeff = 10'sd12; 
			9'd226:  coeff = -10'sd11; 
			9'd227:  coeff = 10'sd9; 
			9'd228:  coeff = -10'sd6; 
			9'd229:  coeff = 10'sd3; 
			9'd230:  coeff = 10'sd0; 
			9'd231:  coeff = -10'sd3; 
			9'd232:  coeff = 10'sd5; 
			9'd233:  coeff = -10'sd7; 
			9'd234:  coeff = 10'sd8; 
			9'd235:  coeff = -10'sd8; 
			9'd236:  coeff = 10'sd7; 
			9'd237:  coeff = -10'sd6; 
			9'd238:  coeff = 10'sd4; 
			9'd239:  coeff = -10'sd2; 
			9'd240:  coeff = 10'sd0; 
			9'd241:  coeff = 10'sd2; 
			9'd242:  coeff = -10'sd4; 
			9'd243:  coeff = 10'sd5; 
			9'd244:  coeff = -10'sd5; 
			9'd245:  coeff = 10'sd6; 
			9'd246:  coeff = -10'sd5; 
			9'd247:  coeff = 10'sd4; 
			9'd248:  coeff = -10'sd3; 
			9'd249:  coeff = 10'sd1; 
			9'd250:  coeff = 10'sd0; 
			9'd251:  coeff = -10'sd1; 
			9'd252:  coeff = 10'sd3; 
			9'd253:  coeff = -10'sd3; 
			9'd254:  coeff = 10'sd4; 
			9'd255:  coeff = -10'sd4; 
			9'd256:  coeff = 10'sd4; 
			9'd257:  coeff = -10'sd3; 
			9'd258:  coeff = 10'sd2; 
			9'd259:  coeff = -10'sd1; 
			9'd260:  coeff = 10'sd0; 
			9'd261:  coeff = 10'sd1; 
			9'd262:  coeff = -10'sd2; 
			9'd263:  coeff = 10'sd2; 
			9'd264:  coeff = -10'sd3; 
			9'd265:  coeff = 10'sd3; 
			9'd266:  coeff = -10'sd3; 
			9'd267:  coeff = 10'sd2; 
			9'd268:  coeff = -10'sd1; 
			9'd269:  coeff = 10'sd1; 
			9'd270:  coeff = 10'sd0; 
			9'd271:  coeff = -10'sd1; 
			9'd272:  coeff = 10'sd1; 
			9'd273:  coeff = -10'sd2; 
			9'd274:  coeff = 10'sd2; 
			9'd275:  coeff = -10'sd2; 
			9'd276:  coeff = 10'sd2; 
			9'd277:  coeff = -10'sd2; 
			9'd278:  coeff = 10'sd1; 
			9'd279:  coeff = -10'sd1; 
			9'd280:  coeff = 10'sd0; 
			9'd281:  coeff = 10'sd0; 
			9'd282:  coeff = -10'sd1; 
			9'd283:  coeff = 10'sd1; 
			9'd284:  coeff = -10'sd1; 
			9'd285:  coeff = 10'sd1; 
			9'd286:  coeff = -10'sd1; 
			9'd287:  coeff = 10'sd1; 
			9'd288:  coeff = -10'sd1; 
			9'd289:  coeff = 10'sd0; 
			9'd290:  coeff = 10'sd0; 
			9'd291:  coeff = 10'sd0; 
			9'd292:  coeff = 10'sd1; 
			9'd293:  coeff = -10'sd1; 
			9'd294:  coeff = 10'sd1; 
			9'd295:  coeff = -10'sd1; 
			9'd296:  coeff = 10'sd1; 
			9'd297:  coeff = -10'sd1; 
			9'd298:  coeff = 10'sd0; 
			9'd299:  coeff = 10'sd0; 
			9'd300:  coeff = 10'sd0; 
			9'd301:  coeff = 10'sd0; 
			9'd302:  coeff = 10'sd0; 
			9'd303:  coeff = 10'sd1; 
			9'd304:  coeff = -10'sd1; 
			9'd305:  coeff = 10'sd1; 
			9'd306:  coeff = -10'sd1; 
			9'd307:  coeff = 10'sd0; 
			9'd308:  coeff = 10'sd0; 
			9'd309:  coeff = 10'sd0; 
			9'd310:  coeff = 10'sd0; 
			9'd311:  coeff = 10'sd0; 
			9'd312:  coeff = 10'sd0; 
			9'd313:  coeff = 10'sd0; 
			9'd314:  coeff = 10'sd0; 
			9'd315:  coeff = 10'sd0; 
			9'd316:  coeff = 10'sd0; 
			9'd317:  coeff = 10'sd0; 
			9'd318:  coeff = 10'sd0; 
			9'd319:  coeff = 10'sd0; 
			9'd320:  coeff = 10'sd0; 
			9'd321:  coeff = 10'sd0; 
			9'd322:  coeff = 10'sd0; 
			9'd323:  coeff = 10'sd0; 
			9'd324:  coeff = 10'sd0; 
			9'd325:  coeff = 10'sd0; 
			9'd326:  coeff = 10'sd0; 
			9'd327:  coeff = 10'sd0; 
			9'd328:  coeff = 10'sd0; 
			9'd329:  coeff = 10'sd0; 
			9'd330:  coeff = 10'sd0; 
			9'd331:  coeff = 10'sd0; 
			9'd332:  coeff = 10'sd0; 
			9'd333:  coeff = 10'sd0; 
			9'd334:  coeff = 10'sd0; 
			9'd335:  coeff = 10'sd0; 
			9'd336:  coeff = 10'sd0; 
			9'd337:  coeff = 10'sd0; 
			9'd338:  coeff = 10'sd0; 
			9'd339:  coeff = 10'sd0; 
			9'd340:  coeff = 10'sd0; 
			9'd341:  coeff = 10'sd0; 
			9'd342:  coeff = 10'sd0; 
			9'd343:  coeff = 10'sd0; 
			9'd344:  coeff = 10'sd0; 
			9'd345:  coeff = 10'sd0; 
			9'd346:  coeff = 10'sd0; 
			9'd347:  coeff = 10'sd0; 
			9'd348:  coeff = 10'sd0; 
			9'd349:  coeff = 10'sd0; 
			9'd350:  coeff = 10'sd0; 
			9'd351:  coeff = 10'sd0; 
			9'd352:  coeff = 10'sd0; 
			9'd353:  coeff = 10'sd0; 
			9'd354:  coeff = 10'sd0; 
			9'd355:  coeff = 10'sd0; 
			9'd356:  coeff = 10'sd0; 
			9'd357:  coeff = 10'sd0; 
			9'd358:  coeff = 10'sd0; 
			9'd359:  coeff = 10'sd0; 
			9'd360:  coeff = 10'sd0; 
			9'd361:  coeff = 10'sd0; 
			9'd362:  coeff = 10'sd0; 
			9'd363:  coeff = 10'sd0; 
			9'd364:  coeff = 10'sd0; 
			9'd365:  coeff = 10'sd0; 
			9'd366:  coeff = 10'sd0; 
			9'd367:  coeff = 10'sd0; 
			9'd368:  coeff = 10'sd0; 
			9'd369:  coeff = 10'sd0; 
			9'd370:  coeff = 10'sd0; 
			9'd371:  coeff = 10'sd0; 
			9'd372:  coeff = 10'sd0; 
			9'd373:  coeff = 10'sd0; 
			9'd374:  coeff = 10'sd0; 
			9'd375:  coeff = 10'sd0; 
			9'd376:  coeff = 10'sd0; 
			9'd377:  coeff = 10'sd0; 
			9'd378:  coeff = 10'sd0; 
			9'd379:  coeff = 10'sd0; 
			9'd380:  coeff = 10'sd0; 
			9'd381:  coeff = 10'sd0; 
			9'd382:  coeff = 10'sd0; 
			9'd383:  coeff = 10'sd0; 
			9'd384:  coeff = 10'sd0; 
			9'd385:  coeff = 10'sd0; 
			9'd386:  coeff = 10'sd0; 
			9'd387:  coeff = 10'sd0; 
			9'd388:  coeff = 10'sd0; 
			9'd389:  coeff = 10'sd0; 
			9'd390:  coeff = 10'sd0; 
			9'd391:  coeff = 10'sd0; 
			9'd392:  coeff = 10'sd0; 
			9'd393:  coeff = 10'sd0; 
			9'd394:  coeff = 10'sd0; 
			9'd395:  coeff = 10'sd0; 
			9'd396:  coeff = 10'sd0; 
			9'd397:  coeff = 10'sd0; 
			9'd398:  coeff = 10'sd0; 
			9'd399:  coeff = 10'sd0; 
			9'd400:  coeff = 10'sd0; 

			default: coeff = 10'hXXX;
		endcase
endmodule

module coeffs400tap_120_260Hz(
  input wire [8:0] index,
  output reg signed [9:0] coeff
);
  // tools will turn this into a 400x10 ROM
	always @(index)
		case (index)
		
			9'd0:  coeff = 10'sd0; 
			9'd1:  coeff = 10'sd0; 
			9'd2:  coeff = 10'sd0; 
			9'd3:  coeff = 10'sd0; 
			9'd4:  coeff = 10'sd0; 
			9'd5:  coeff = 10'sd0; 
			9'd6:  coeff = 10'sd0; 
			9'd7:  coeff = 10'sd0; 
			9'd8:  coeff = 10'sd0; 
			9'd9:  coeff = 10'sd0; 
			9'd10:  coeff = 10'sd0; 
			9'd11:  coeff = 10'sd0; 
			9'd12:  coeff = 10'sd0; 
			9'd13:  coeff = 10'sd0; 
			9'd14:  coeff = 10'sd0; 
			9'd15:  coeff = 10'sd0; 
			9'd16:  coeff = 10'sd0; 
			9'd17:  coeff = 10'sd0; 
			9'd18:  coeff = 10'sd0; 
			9'd19:  coeff = 10'sd0; 
			9'd20:  coeff = 10'sd0; 
			9'd21:  coeff = 10'sd0; 
			9'd22:  coeff = 10'sd0; 
			9'd23:  coeff = 10'sd0; 
			9'd24:  coeff = 10'sd0; 
			9'd25:  coeff = 10'sd0; 
			9'd26:  coeff = 10'sd0; 
			9'd27:  coeff = 10'sd0; 
			9'd28:  coeff = 10'sd0; 
			9'd29:  coeff = 10'sd0; 
			9'd30:  coeff = 10'sd0; 
			9'd31:  coeff = 10'sd0; 
			9'd32:  coeff = 10'sd0; 
			9'd33:  coeff = 10'sd0; 
			9'd34:  coeff = 10'sd0; 
			9'd35:  coeff = 10'sd0; 
			9'd36:  coeff = 10'sd0; 
			9'd37:  coeff = 10'sd0; 
			9'd38:  coeff = 10'sd0; 
			9'd39:  coeff = 10'sd0; 
			9'd40:  coeff = 10'sd0; 
			9'd41:  coeff = 10'sd0; 
			9'd42:  coeff = 10'sd0; 
			9'd43:  coeff = 10'sd0; 
			9'd44:  coeff = 10'sd0; 
			9'd45:  coeff = 10'sd0; 
			9'd46:  coeff = 10'sd0; 
			9'd47:  coeff = 10'sd0; 
			9'd48:  coeff = 10'sd0; 
			9'd49:  coeff = 10'sd0; 
			9'd50:  coeff = 10'sd0; 
			9'd51:  coeff = 10'sd0; 
			9'd52:  coeff = 10'sd0; 
			9'd53:  coeff = 10'sd0; 
			9'd54:  coeff = 10'sd0; 
			9'd55:  coeff = 10'sd0; 
			9'd56:  coeff = 10'sd0; 
			9'd57:  coeff = 10'sd0; 
			9'd58:  coeff = 10'sd0; 
			9'd59:  coeff = 10'sd0; 
			9'd60:  coeff = 10'sd0; 
			9'd61:  coeff = -10'sd1; 
			9'd62:  coeff = -10'sd1; 
			9'd63:  coeff = -10'sd1; 
			9'd64:  coeff = -10'sd1; 
			9'd65:  coeff = -10'sd1; 
			9'd66:  coeff = -10'sd1; 
			9'd67:  coeff = -10'sd1; 
			9'd68:  coeff = -10'sd1; 
			9'd69:  coeff = -10'sd1; 
			9'd70:  coeff = -10'sd1; 
			9'd71:  coeff = -10'sd1; 
			9'd72:  coeff = -10'sd1; 
			9'd73:  coeff = -10'sd1; 
			9'd74:  coeff = -10'sd1; 
			9'd75:  coeff = -10'sd1; 
			9'd76:  coeff = -10'sd1; 
			9'd77:  coeff = -10'sd1; 
			9'd78:  coeff = -10'sd1; 
			9'd79:  coeff = -10'sd1; 
			9'd80:  coeff = -10'sd1; 
			9'd81:  coeff = -10'sd1; 
			9'd82:  coeff = -10'sd1; 
			9'd83:  coeff = -10'sd2; 
			9'd84:  coeff = -10'sd2; 
			9'd85:  coeff = -10'sd2; 
			9'd86:  coeff = -10'sd2; 
			9'd87:  coeff = -10'sd2; 
			9'd88:  coeff = -10'sd2; 
			9'd89:  coeff = -10'sd2; 
			9'd90:  coeff = -10'sd2; 
			9'd91:  coeff = -10'sd2; 
			9'd92:  coeff = -10'sd2; 
			9'd93:  coeff = -10'sd2; 
			9'd94:  coeff = -10'sd2; 
			9'd95:  coeff = -10'sd2; 
			9'd96:  coeff = -10'sd2; 
			9'd97:  coeff = -10'sd2; 
			9'd98:  coeff = -10'sd2; 
			9'd99:  coeff = -10'sd2; 
			9'd100:  coeff = -10'sd2; 
			9'd101:  coeff = -10'sd2; 
			9'd102:  coeff = -10'sd2; 
			9'd103:  coeff = -10'sd2; 
			9'd104:  coeff = -10'sd3; 
			9'd105:  coeff = -10'sd3; 
			9'd106:  coeff = -10'sd3; 
			9'd107:  coeff = -10'sd3; 
			9'd108:  coeff = -10'sd3; 
			9'd109:  coeff = -10'sd3; 
			9'd110:  coeff = -10'sd3; 
			9'd111:  coeff = -10'sd3; 
			9'd112:  coeff = -10'sd3; 
			9'd113:  coeff = -10'sd3; 
			9'd114:  coeff = -10'sd3; 
			9'd115:  coeff = -10'sd3; 
			9'd116:  coeff = -10'sd2; 
			9'd117:  coeff = -10'sd2; 
			9'd118:  coeff = -10'sd2; 
			9'd119:  coeff = -10'sd2; 
			9'd120:  coeff = -10'sd2; 
			9'd121:  coeff = -10'sd2; 
			9'd122:  coeff = -10'sd2; 
			9'd123:  coeff = -10'sd2; 
			9'd124:  coeff = -10'sd2; 
			9'd125:  coeff = -10'sd2; 
			9'd126:  coeff = -10'sd2; 
			9'd127:  coeff = -10'sd2; 
			9'd128:  coeff = -10'sd2; 
			9'd129:  coeff = -10'sd1; 
			9'd130:  coeff = -10'sd1; 
			9'd131:  coeff = -10'sd1; 
			9'd132:  coeff = -10'sd1; 
			9'd133:  coeff = -10'sd1; 
			9'd134:  coeff = -10'sd1; 
			9'd135:  coeff = 10'sd0; 
			9'd136:  coeff = 10'sd0; 
			9'd137:  coeff = 10'sd0; 
			9'd138:  coeff = 10'sd0; 
			9'd139:  coeff = 10'sd0; 
			9'd140:  coeff = 10'sd1; 
			9'd141:  coeff = 10'sd1; 
			9'd142:  coeff = 10'sd1; 
			9'd143:  coeff = 10'sd1; 
			9'd144:  coeff = 10'sd1; 
			9'd145:  coeff = 10'sd2; 
			9'd146:  coeff = 10'sd2; 
			9'd147:  coeff = 10'sd2; 
			9'd148:  coeff = 10'sd2; 
			9'd149:  coeff = 10'sd3; 
			9'd150:  coeff = 10'sd3; 
			9'd151:  coeff = 10'sd3; 
			9'd152:  coeff = 10'sd4; 
			9'd153:  coeff = 10'sd4; 
			9'd154:  coeff = 10'sd4; 
			9'd155:  coeff = 10'sd5; 
			9'd156:  coeff = 10'sd5; 
			9'd157:  coeff = 10'sd5; 
			9'd158:  coeff = 10'sd5; 
			9'd159:  coeff = 10'sd6; 
			9'd160:  coeff = 10'sd6; 
			9'd161:  coeff = 10'sd6; 
			9'd162:  coeff = 10'sd7; 
			9'd163:  coeff = 10'sd7; 
			9'd164:  coeff = 10'sd7; 
			9'd165:  coeff = 10'sd8; 
			9'd166:  coeff = 10'sd8; 
			9'd167:  coeff = 10'sd8; 
			9'd168:  coeff = 10'sd9; 
			9'd169:  coeff = 10'sd9; 
			9'd170:  coeff = 10'sd9; 
			9'd171:  coeff = 10'sd9; 
			9'd172:  coeff = 10'sd10; 
			9'd173:  coeff = 10'sd10; 
			9'd174:  coeff = 10'sd10; 
			9'd175:  coeff = 10'sd11; 
			9'd176:  coeff = 10'sd11; 
			9'd177:  coeff = 10'sd11; 
			9'd178:  coeff = 10'sd11; 
			9'd179:  coeff = 10'sd12; 
			9'd180:  coeff = 10'sd12; 
			9'd181:  coeff = 10'sd12; 
			9'd182:  coeff = 10'sd12; 
			9'd183:  coeff = 10'sd12; 
			9'd184:  coeff = 10'sd13; 
			9'd185:  coeff = 10'sd13; 
			9'd186:  coeff = 10'sd13; 
			9'd187:  coeff = 10'sd13; 
			9'd188:  coeff = 10'sd13; 
			9'd189:  coeff = 10'sd14; 
			9'd190:  coeff = 10'sd14; 
			9'd191:  coeff = 10'sd14; 
			9'd192:  coeff = 10'sd14; 
			9'd193:  coeff = 10'sd14; 
			9'd194:  coeff = 10'sd14; 
			9'd195:  coeff = 10'sd14; 
			9'd196:  coeff = 10'sd14; 
			9'd197:  coeff = 10'sd14; 
			9'd198:  coeff = 10'sd14; 
			9'd199:  coeff = 10'sd14; 
			9'd200:  coeff = 10'sd14; 
			9'd201:  coeff = 10'sd14; 
			9'd202:  coeff = 10'sd14; 
			9'd203:  coeff = 10'sd14; 
			9'd204:  coeff = 10'sd14; 
			9'd205:  coeff = 10'sd14; 
			9'd206:  coeff = 10'sd14; 
			9'd207:  coeff = 10'sd14; 
			9'd208:  coeff = 10'sd14; 
			9'd209:  coeff = 10'sd14; 
			9'd210:  coeff = 10'sd14; 
			9'd211:  coeff = 10'sd14; 
			9'd212:  coeff = 10'sd13; 
			9'd213:  coeff = 10'sd13; 
			9'd214:  coeff = 10'sd13; 
			9'd215:  coeff = 10'sd13; 
			9'd216:  coeff = 10'sd13; 
			9'd217:  coeff = 10'sd12; 
			9'd218:  coeff = 10'sd12; 
			9'd219:  coeff = 10'sd12; 
			9'd220:  coeff = 10'sd12; 
			9'd221:  coeff = 10'sd12; 
			9'd222:  coeff = 10'sd11; 
			9'd223:  coeff = 10'sd11; 
			9'd224:  coeff = 10'sd11; 
			9'd225:  coeff = 10'sd11; 
			9'd226:  coeff = 10'sd10; 
			9'd227:  coeff = 10'sd10; 
			9'd228:  coeff = 10'sd10; 
			9'd229:  coeff = 10'sd9; 
			9'd230:  coeff = 10'sd9; 
			9'd231:  coeff = 10'sd9; 
			9'd232:  coeff = 10'sd9; 
			9'd233:  coeff = 10'sd8; 
			9'd234:  coeff = 10'sd8; 
			9'd235:  coeff = 10'sd8; 
			9'd236:  coeff = 10'sd7; 
			9'd237:  coeff = 10'sd7; 
			9'd238:  coeff = 10'sd7; 
			9'd239:  coeff = 10'sd6; 
			9'd240:  coeff = 10'sd6; 
			9'd241:  coeff = 10'sd6; 
			9'd242:  coeff = 10'sd5; 
			9'd243:  coeff = 10'sd5; 
			9'd244:  coeff = 10'sd5; 
			9'd245:  coeff = 10'sd5; 
			9'd246:  coeff = 10'sd4; 
			9'd247:  coeff = 10'sd4; 
			9'd248:  coeff = 10'sd4; 
			9'd249:  coeff = 10'sd3; 
			9'd250:  coeff = 10'sd3; 
			9'd251:  coeff = 10'sd3; 
			9'd252:  coeff = 10'sd2; 
			9'd253:  coeff = 10'sd2; 
			9'd254:  coeff = 10'sd2; 
			9'd255:  coeff = 10'sd2; 
			9'd256:  coeff = 10'sd1; 
			9'd257:  coeff = 10'sd1; 
			9'd258:  coeff = 10'sd1; 
			9'd259:  coeff = 10'sd1; 
			9'd260:  coeff = 10'sd1; 
			9'd261:  coeff = 10'sd0; 
			9'd262:  coeff = 10'sd0; 
			9'd263:  coeff = 10'sd0; 
			9'd264:  coeff = 10'sd0; 
			9'd265:  coeff = 10'sd0; 
			9'd266:  coeff = -10'sd1; 
			9'd267:  coeff = -10'sd1; 
			9'd268:  coeff = -10'sd1; 
			9'd269:  coeff = -10'sd1; 
			9'd270:  coeff = -10'sd1; 
			9'd271:  coeff = -10'sd1; 
			9'd272:  coeff = -10'sd2; 
			9'd273:  coeff = -10'sd2; 
			9'd274:  coeff = -10'sd2; 
			9'd275:  coeff = -10'sd2; 
			9'd276:  coeff = -10'sd2; 
			9'd277:  coeff = -10'sd2; 
			9'd278:  coeff = -10'sd2; 
			9'd279:  coeff = -10'sd2; 
			9'd280:  coeff = -10'sd2; 
			9'd281:  coeff = -10'sd2; 
			9'd282:  coeff = -10'sd2; 
			9'd283:  coeff = -10'sd2; 
			9'd284:  coeff = -10'sd2; 
			9'd285:  coeff = -10'sd3; 
			9'd286:  coeff = -10'sd3; 
			9'd287:  coeff = -10'sd3; 
			9'd288:  coeff = -10'sd3; 
			9'd289:  coeff = -10'sd3; 
			9'd290:  coeff = -10'sd3; 
			9'd291:  coeff = -10'sd3; 
			9'd292:  coeff = -10'sd3; 
			9'd293:  coeff = -10'sd3; 
			9'd294:  coeff = -10'sd3; 
			9'd295:  coeff = -10'sd3; 
			9'd296:  coeff = -10'sd3; 
			9'd297:  coeff = -10'sd2; 
			9'd298:  coeff = -10'sd2; 
			9'd299:  coeff = -10'sd2; 
			9'd300:  coeff = -10'sd2; 
			9'd301:  coeff = -10'sd2; 
			9'd302:  coeff = -10'sd2; 
			9'd303:  coeff = -10'sd2; 
			9'd304:  coeff = -10'sd2; 
			9'd305:  coeff = -10'sd2; 
			9'd306:  coeff = -10'sd2; 
			9'd307:  coeff = -10'sd2; 
			9'd308:  coeff = -10'sd2; 
			9'd309:  coeff = -10'sd2; 
			9'd310:  coeff = -10'sd2; 
			9'd311:  coeff = -10'sd2; 
			9'd312:  coeff = -10'sd2; 
			9'd313:  coeff = -10'sd2; 
			9'd314:  coeff = -10'sd2; 
			9'd315:  coeff = -10'sd2; 
			9'd316:  coeff = -10'sd2; 
			9'd317:  coeff = -10'sd2; 
			9'd318:  coeff = -10'sd1; 
			9'd319:  coeff = -10'sd1; 
			9'd320:  coeff = -10'sd1; 
			9'd321:  coeff = -10'sd1; 
			9'd322:  coeff = -10'sd1; 
			9'd323:  coeff = -10'sd1; 
			9'd324:  coeff = -10'sd1; 
			9'd325:  coeff = -10'sd1; 
			9'd326:  coeff = -10'sd1; 
			9'd327:  coeff = -10'sd1; 
			9'd328:  coeff = -10'sd1; 
			9'd329:  coeff = -10'sd1; 
			9'd330:  coeff = -10'sd1; 
			9'd331:  coeff = -10'sd1; 
			9'd332:  coeff = -10'sd1; 
			9'd333:  coeff = -10'sd1; 
			9'd334:  coeff = -10'sd1; 
			9'd335:  coeff = -10'sd1; 
			9'd336:  coeff = -10'sd1; 
			9'd337:  coeff = -10'sd1; 
			9'd338:  coeff = -10'sd1; 
			9'd339:  coeff = -10'sd1; 
			9'd340:  coeff = 10'sd0; 
			9'd341:  coeff = 10'sd0; 
			9'd342:  coeff = 10'sd0; 
			9'd343:  coeff = 10'sd0; 
			9'd344:  coeff = 10'sd0; 
			9'd345:  coeff = 10'sd0; 
			9'd346:  coeff = 10'sd0; 
			9'd347:  coeff = 10'sd0; 
			9'd348:  coeff = 10'sd0; 
			9'd349:  coeff = 10'sd0; 
			9'd350:  coeff = 10'sd0; 
			9'd351:  coeff = 10'sd0; 
			9'd352:  coeff = 10'sd0; 
			9'd353:  coeff = 10'sd0; 
			9'd354:  coeff = 10'sd0; 
			9'd355:  coeff = 10'sd0; 
			9'd356:  coeff = 10'sd0; 
			9'd357:  coeff = 10'sd0; 
			9'd358:  coeff = 10'sd0; 
			9'd359:  coeff = 10'sd0; 
			9'd360:  coeff = 10'sd0; 
			9'd361:  coeff = 10'sd0; 
			9'd362:  coeff = 10'sd0; 
			9'd363:  coeff = 10'sd0; 
			9'd364:  coeff = 10'sd0; 
			9'd365:  coeff = 10'sd0; 
			9'd366:  coeff = 10'sd0; 
			9'd367:  coeff = 10'sd0; 
			9'd368:  coeff = 10'sd0; 
			9'd369:  coeff = 10'sd0; 
			9'd370:  coeff = 10'sd0; 
			9'd371:  coeff = 10'sd0; 
			9'd372:  coeff = 10'sd0; 
			9'd373:  coeff = 10'sd0; 
			9'd374:  coeff = 10'sd0; 
			9'd375:  coeff = 10'sd0; 
			9'd376:  coeff = 10'sd0; 
			9'd377:  coeff = 10'sd0; 
			9'd378:  coeff = 10'sd0; 
			9'd379:  coeff = 10'sd0; 
			9'd380:  coeff = 10'sd0; 
			9'd381:  coeff = 10'sd0; 
			9'd382:  coeff = 10'sd0; 
			9'd383:  coeff = 10'sd0; 
			9'd384:  coeff = 10'sd0; 
			9'd385:  coeff = 10'sd0; 
			9'd386:  coeff = 10'sd0; 
			9'd387:  coeff = 10'sd0; 
			9'd388:  coeff = 10'sd0; 
			9'd389:  coeff = 10'sd0; 
			9'd390:  coeff = 10'sd0; 
			9'd391:  coeff = 10'sd0; 
			9'd392:  coeff = 10'sd0; 
			9'd393:  coeff = 10'sd0; 
			9'd394:  coeff = 10'sd0; 
			9'd395:  coeff = 10'sd0; 
			9'd396:  coeff = 10'sd0; 
			9'd397:  coeff = 10'sd0; 
			9'd398:  coeff = 10'sd0; 
			9'd399:  coeff = 10'sd0; 
			9'd400:  coeff = 10'sd0; 

			default: coeff = 10'hXXX;
		endcase
endmodule

module coeffs400tap_260_600Hz(
  input wire [8:0] index,
  output reg signed [9:0] coeff
);
  // tools will turn this into a 401x10 ROM
	always @(index)
		case (index)

			9'd0:  coeff = 10'sd0; 
			9'd1:  coeff = 10'sd0; 
			9'd2:  coeff = 10'sd0; 
			9'd3:  coeff = 10'sd0; 
			9'd4:  coeff = 10'sd0; 
			9'd5:  coeff = 10'sd0; 
			9'd6:  coeff = 10'sd0; 
			9'd7:  coeff = 10'sd0; 
			9'd8:  coeff = 10'sd0; 
			9'd9:  coeff = 10'sd0; 
			9'd10:  coeff = 10'sd0; 
			9'd11:  coeff = 10'sd0; 
			9'd12:  coeff = 10'sd0; 
			9'd13:  coeff = 10'sd0; 
			9'd14:  coeff = 10'sd0; 
			9'd15:  coeff = 10'sd0; 
			9'd16:  coeff = 10'sd0; 
			9'd17:  coeff = 10'sd0; 
			9'd18:  coeff = 10'sd0; 
			9'd19:  coeff = 10'sd0; 
			9'd20:  coeff = 10'sd0; 
			9'd21:  coeff = 10'sd0; 
			9'd22:  coeff = 10'sd0; 
			9'd23:  coeff = 10'sd0; 
			9'd24:  coeff = 10'sd0; 
			9'd25:  coeff = 10'sd0; 
			9'd26:  coeff = 10'sd0; 
			9'd27:  coeff = 10'sd0; 
			9'd28:  coeff = 10'sd0; 
			9'd29:  coeff = 10'sd0; 
			9'd30:  coeff = 10'sd0; 
			9'd31:  coeff = 10'sd0; 
			9'd32:  coeff = 10'sd0; 
			9'd33:  coeff = 10'sd0; 
			9'd34:  coeff = 10'sd0; 
			9'd35:  coeff = 10'sd0; 
			9'd36:  coeff = 10'sd0; 
			9'd37:  coeff = 10'sd0; 
			9'd38:  coeff = 10'sd0; 
			9'd39:  coeff = 10'sd0; 
			9'd40:  coeff = 10'sd0; 
			9'd41:  coeff = 10'sd0; 
			9'd42:  coeff = 10'sd0; 
			9'd43:  coeff = 10'sd0; 
			9'd44:  coeff = 10'sd0; 
			9'd45:  coeff = 10'sd0; 
			9'd46:  coeff = 10'sd0; 
			9'd47:  coeff = 10'sd0; 
			9'd48:  coeff = 10'sd0; 
			9'd49:  coeff = 10'sd0; 
			9'd50:  coeff = 10'sd0; 
			9'd51:  coeff = 10'sd0; 
			9'd52:  coeff = 10'sd0; 
			9'd53:  coeff = 10'sd0; 
			9'd54:  coeff = 10'sd0; 
			9'd55:  coeff = 10'sd0; 
			9'd56:  coeff = 10'sd0; 
			9'd57:  coeff = 10'sd0; 
			9'd58:  coeff = 10'sd0; 
			9'd59:  coeff = 10'sd0; 
			9'd60:  coeff = 10'sd0; 
			9'd61:  coeff = 10'sd0; 
			9'd62:  coeff = 10'sd0; 
			9'd63:  coeff = 10'sd0; 
			9'd64:  coeff = 10'sd0; 
			9'd65:  coeff = 10'sd0; 
			9'd66:  coeff = 10'sd0; 
			9'd67:  coeff = 10'sd0; 
			9'd68:  coeff = 10'sd0; 
			9'd69:  coeff = 10'sd0; 
			9'd70:  coeff = 10'sd0; 
			9'd71:  coeff = 10'sd0; 
			9'd72:  coeff = 10'sd0; 
			9'd73:  coeff = 10'sd0; 
			9'd74:  coeff = 10'sd0; 
			9'd75:  coeff = 10'sd0; 
			9'd76:  coeff = 10'sd0; 
			9'd77:  coeff = 10'sd0; 
			9'd78:  coeff = 10'sd0; 
			9'd79:  coeff = 10'sd0; 
			9'd80:  coeff = 10'sd0; 
			9'd81:  coeff = 10'sd0; 
			9'd82:  coeff = 10'sd0; 
			9'd83:  coeff = 10'sd0; 
			9'd84:  coeff = 10'sd1; 
			9'd85:  coeff = 10'sd1; 
			9'd86:  coeff = 10'sd1; 
			9'd87:  coeff = 10'sd1; 
			9'd88:  coeff = 10'sd1; 
			9'd89:  coeff = 10'sd1; 
			9'd90:  coeff = 10'sd1; 
			9'd91:  coeff = 10'sd1; 
			9'd92:  coeff = 10'sd1; 
			9'd93:  coeff = 10'sd1; 
			9'd94:  coeff = 10'sd1; 
			9'd95:  coeff = 10'sd1; 
			9'd96:  coeff = 10'sd1; 
			9'd97:  coeff = 10'sd1; 
			9'd98:  coeff = 10'sd1; 
			9'd99:  coeff = 10'sd1; 
			9'd100:  coeff = 10'sd1; 
			9'd101:  coeff = 10'sd1; 
			9'd102:  coeff = 10'sd1; 
			9'd103:  coeff = 10'sd1; 
			9'd104:  coeff = 10'sd1; 
			9'd105:  coeff = 10'sd1; 
			9'd106:  coeff = 10'sd1; 
			9'd107:  coeff = 10'sd1; 
			9'd108:  coeff = 10'sd1; 
			9'd109:  coeff = 10'sd1; 
			9'd110:  coeff = 10'sd1; 
			9'd111:  coeff = 10'sd1; 
			9'd112:  coeff = 10'sd1; 
			9'd113:  coeff = 10'sd1; 
			9'd114:  coeff = 10'sd0; 
			9'd115:  coeff = 10'sd0; 
			9'd116:  coeff = 10'sd0; 
			9'd117:  coeff = 10'sd0; 
			9'd118:  coeff = 10'sd0; 
			9'd119:  coeff = -10'sd1; 
			9'd120:  coeff = -10'sd1; 
			9'd121:  coeff = -10'sd1; 
			9'd122:  coeff = -10'sd1; 
			9'd123:  coeff = -10'sd2; 
			9'd124:  coeff = -10'sd2; 
			9'd125:  coeff = -10'sd2; 
			9'd126:  coeff = -10'sd3; 
			9'd127:  coeff = -10'sd3; 
			9'd128:  coeff = -10'sd3; 
			9'd129:  coeff = -10'sd4; 
			9'd130:  coeff = -10'sd4; 
			9'd131:  coeff = -10'sd4; 
			9'd132:  coeff = -10'sd5; 
			9'd133:  coeff = -10'sd5; 
			9'd134:  coeff = -10'sd5; 
			9'd135:  coeff = -10'sd6; 
			9'd136:  coeff = -10'sd6; 
			9'd137:  coeff = -10'sd7; 
			9'd138:  coeff = -10'sd7; 
			9'd139:  coeff = -10'sd7; 
			9'd140:  coeff = -10'sd8; 
			9'd141:  coeff = -10'sd8; 
			9'd142:  coeff = -10'sd8; 
			9'd143:  coeff = -10'sd9; 
			9'd144:  coeff = -10'sd9; 
			9'd145:  coeff = -10'sd9; 
			9'd146:  coeff = -10'sd9; 
			9'd147:  coeff = -10'sd9; 
			9'd148:  coeff = -10'sd9; 
			9'd149:  coeff = -10'sd10; 
			9'd150:  coeff = -10'sd10; 
			9'd151:  coeff = -10'sd10; 
			9'd152:  coeff = -10'sd10; 
			9'd153:  coeff = -10'sd10; 
			9'd154:  coeff = -10'sd9; 
			9'd155:  coeff = -10'sd9; 
			9'd156:  coeff = -10'sd9; 
			9'd157:  coeff = -10'sd9; 
			9'd158:  coeff = -10'sd9; 
			9'd159:  coeff = -10'sd8; 
			9'd160:  coeff = -10'sd8; 
			9'd161:  coeff = -10'sd7; 
			9'd162:  coeff = -10'sd7; 
			9'd163:  coeff = -10'sd7; 
			9'd164:  coeff = -10'sd6; 
			9'd165:  coeff = -10'sd5; 
			9'd166:  coeff = -10'sd5; 
			9'd167:  coeff = -10'sd4; 
			9'd168:  coeff = -10'sd3; 
			9'd169:  coeff = -10'sd3; 
			9'd170:  coeff = -10'sd2; 
			9'd171:  coeff = -10'sd1; 
			9'd172:  coeff = 10'sd0; 
			9'd173:  coeff = 10'sd1; 
			9'd174:  coeff = 10'sd2; 
			9'd175:  coeff = 10'sd2; 
			9'd176:  coeff = 10'sd3; 
			9'd177:  coeff = 10'sd4; 
			9'd178:  coeff = 10'sd5; 
			9'd179:  coeff = 10'sd6; 
			9'd180:  coeff = 10'sd7; 
			9'd181:  coeff = 10'sd8; 
			9'd182:  coeff = 10'sd9; 
			9'd183:  coeff = 10'sd9; 
			9'd184:  coeff = 10'sd10; 
			9'd185:  coeff = 10'sd11; 
			9'd186:  coeff = 10'sd12; 
			9'd187:  coeff = 10'sd13; 
			9'd188:  coeff = 10'sd13; 
			9'd189:  coeff = 10'sd14; 
			9'd190:  coeff = 10'sd15; 
			9'd191:  coeff = 10'sd15; 
			9'd192:  coeff = 10'sd16; 
			9'd193:  coeff = 10'sd16; 
			9'd194:  coeff = 10'sd16; 
			9'd195:  coeff = 10'sd17; 
			9'd196:  coeff = 10'sd17; 
			9'd197:  coeff = 10'sd17; 
			9'd198:  coeff = 10'sd17; 
			9'd199:  coeff = 10'sd18; 
			9'd200:  coeff = 10'sd18; 
			9'd201:  coeff = 10'sd18; 
			9'd202:  coeff = 10'sd17; 
			9'd203:  coeff = 10'sd17; 
			9'd204:  coeff = 10'sd17; 
			9'd205:  coeff = 10'sd17; 
			9'd206:  coeff = 10'sd16; 
			9'd207:  coeff = 10'sd16; 
			9'd208:  coeff = 10'sd16; 
			9'd209:  coeff = 10'sd15; 
			9'd210:  coeff = 10'sd15; 
			9'd211:  coeff = 10'sd14; 
			9'd212:  coeff = 10'sd13; 
			9'd213:  coeff = 10'sd13; 
			9'd214:  coeff = 10'sd12; 
			9'd215:  coeff = 10'sd11; 
			9'd216:  coeff = 10'sd10; 
			9'd217:  coeff = 10'sd9; 
			9'd218:  coeff = 10'sd9; 
			9'd219:  coeff = 10'sd8; 
			9'd220:  coeff = 10'sd7; 
			9'd221:  coeff = 10'sd6; 
			9'd222:  coeff = 10'sd5; 
			9'd223:  coeff = 10'sd4; 
			9'd224:  coeff = 10'sd3; 
			9'd225:  coeff = 10'sd2; 
			9'd226:  coeff = 10'sd2; 
			9'd227:  coeff = 10'sd1; 
			9'd228:  coeff = 10'sd0; 
			9'd229:  coeff = -10'sd1; 
			9'd230:  coeff = -10'sd2; 
			9'd231:  coeff = -10'sd3; 
			9'd232:  coeff = -10'sd3; 
			9'd233:  coeff = -10'sd4; 
			9'd234:  coeff = -10'sd5; 
			9'd235:  coeff = -10'sd5; 
			9'd236:  coeff = -10'sd6; 
			9'd237:  coeff = -10'sd7; 
			9'd238:  coeff = -10'sd7; 
			9'd239:  coeff = -10'sd7; 
			9'd240:  coeff = -10'sd8; 
			9'd241:  coeff = -10'sd8; 
			9'd242:  coeff = -10'sd9; 
			9'd243:  coeff = -10'sd9; 
			9'd244:  coeff = -10'sd9; 
			9'd245:  coeff = -10'sd9; 
			9'd246:  coeff = -10'sd9; 
			9'd247:  coeff = -10'sd10; 
			9'd248:  coeff = -10'sd10; 
			9'd249:  coeff = -10'sd10; 
			9'd250:  coeff = -10'sd10; 
			9'd251:  coeff = -10'sd10; 
			9'd252:  coeff = -10'sd9; 
			9'd253:  coeff = -10'sd9; 
			9'd254:  coeff = -10'sd9; 
			9'd255:  coeff = -10'sd9; 
			9'd256:  coeff = -10'sd9; 
			9'd257:  coeff = -10'sd9; 
			9'd258:  coeff = -10'sd8; 
			9'd259:  coeff = -10'sd8; 
			9'd260:  coeff = -10'sd8; 
			9'd261:  coeff = -10'sd7; 
			9'd262:  coeff = -10'sd7; 
			9'd263:  coeff = -10'sd7; 
			9'd264:  coeff = -10'sd6; 
			9'd265:  coeff = -10'sd6; 
			9'd266:  coeff = -10'sd5; 
			9'd267:  coeff = -10'sd5; 
			9'd268:  coeff = -10'sd5; 
			9'd269:  coeff = -10'sd4; 
			9'd270:  coeff = -10'sd4; 
			9'd271:  coeff = -10'sd4; 
			9'd272:  coeff = -10'sd3; 
			9'd273:  coeff = -10'sd3; 
			9'd274:  coeff = -10'sd3; 
			9'd275:  coeff = -10'sd2; 
			9'd276:  coeff = -10'sd2; 
			9'd277:  coeff = -10'sd2; 
			9'd278:  coeff = -10'sd1; 
			9'd279:  coeff = -10'sd1; 
			9'd280:  coeff = -10'sd1; 
			9'd281:  coeff = -10'sd1; 
			9'd282:  coeff = 10'sd0; 
			9'd283:  coeff = 10'sd0; 
			9'd284:  coeff = 10'sd0; 
			9'd285:  coeff = 10'sd0; 
			9'd286:  coeff = 10'sd0; 
			9'd287:  coeff = 10'sd1; 
			9'd288:  coeff = 10'sd1; 
			9'd289:  coeff = 10'sd1; 
			9'd290:  coeff = 10'sd1; 
			9'd291:  coeff = 10'sd1; 
			9'd292:  coeff = 10'sd1; 
			9'd293:  coeff = 10'sd1; 
			9'd294:  coeff = 10'sd1; 
			9'd295:  coeff = 10'sd1; 
			9'd296:  coeff = 10'sd1; 
			9'd297:  coeff = 10'sd1; 
			9'd298:  coeff = 10'sd1; 
			9'd299:  coeff = 10'sd1; 
			9'd300:  coeff = 10'sd1; 
			9'd301:  coeff = 10'sd1; 
			9'd302:  coeff = 10'sd1; 
			9'd303:  coeff = 10'sd1; 
			9'd304:  coeff = 10'sd1; 
			9'd305:  coeff = 10'sd1; 
			9'd306:  coeff = 10'sd1; 
			9'd307:  coeff = 10'sd1; 
			9'd308:  coeff = 10'sd1; 
			9'd309:  coeff = 10'sd1; 
			9'd310:  coeff = 10'sd1; 
			9'd311:  coeff = 10'sd1; 
			9'd312:  coeff = 10'sd1; 
			9'd313:  coeff = 10'sd1; 
			9'd314:  coeff = 10'sd1; 
			9'd315:  coeff = 10'sd1; 
			9'd316:  coeff = 10'sd1; 
			9'd317:  coeff = 10'sd0; 
			9'd318:  coeff = 10'sd0; 
			9'd319:  coeff = 10'sd0; 
			9'd320:  coeff = 10'sd0; 
			9'd321:  coeff = 10'sd0; 
			9'd322:  coeff = 10'sd0; 
			9'd323:  coeff = 10'sd0; 
			9'd324:  coeff = 10'sd0; 
			9'd325:  coeff = 10'sd0; 
			9'd326:  coeff = 10'sd0; 
			9'd327:  coeff = 10'sd0; 
			9'd328:  coeff = 10'sd0; 
			9'd329:  coeff = 10'sd0; 
			9'd330:  coeff = 10'sd0; 
			9'd331:  coeff = 10'sd0; 
			9'd332:  coeff = 10'sd0; 
			9'd333:  coeff = 10'sd0; 
			9'd334:  coeff = 10'sd0; 
			9'd335:  coeff = 10'sd0; 
			9'd336:  coeff = 10'sd0; 
			9'd337:  coeff = 10'sd0; 
			9'd338:  coeff = 10'sd0; 
			9'd339:  coeff = 10'sd0; 
			9'd340:  coeff = 10'sd0; 
			9'd341:  coeff = 10'sd0; 
			9'd342:  coeff = 10'sd0; 
			9'd343:  coeff = 10'sd0; 
			9'd344:  coeff = 10'sd0; 
			9'd345:  coeff = 10'sd0; 
			9'd346:  coeff = 10'sd0; 
			9'd347:  coeff = 10'sd0; 
			9'd348:  coeff = 10'sd0; 
			9'd349:  coeff = 10'sd0; 
			9'd350:  coeff = 10'sd0; 
			9'd351:  coeff = 10'sd0; 
			9'd352:  coeff = 10'sd0; 
			9'd353:  coeff = 10'sd0; 
			9'd354:  coeff = 10'sd0; 
			9'd355:  coeff = 10'sd0; 
			9'd356:  coeff = 10'sd0; 
			9'd357:  coeff = 10'sd0; 
			9'd358:  coeff = 10'sd0; 
			9'd359:  coeff = 10'sd0; 
			9'd360:  coeff = 10'sd0; 
			9'd361:  coeff = 10'sd0; 
			9'd362:  coeff = 10'sd0; 
			9'd363:  coeff = 10'sd0; 
			9'd364:  coeff = 10'sd0; 
			9'd365:  coeff = 10'sd0; 
			9'd366:  coeff = 10'sd0; 
			9'd367:  coeff = 10'sd0; 
			9'd368:  coeff = 10'sd0; 
			9'd369:  coeff = 10'sd0; 
			9'd370:  coeff = 10'sd0; 
			9'd371:  coeff = 10'sd0; 
			9'd372:  coeff = 10'sd0; 
			9'd373:  coeff = 10'sd0; 
			9'd374:  coeff = 10'sd0; 
			9'd375:  coeff = 10'sd0; 
			9'd376:  coeff = 10'sd0; 
			9'd377:  coeff = 10'sd0; 
			9'd378:  coeff = 10'sd0; 
			9'd379:  coeff = 10'sd0; 
			9'd380:  coeff = 10'sd0; 
			9'd381:  coeff = 10'sd0; 
			9'd382:  coeff = 10'sd0; 
			9'd383:  coeff = 10'sd0; 
			9'd384:  coeff = 10'sd0; 
			9'd385:  coeff = 10'sd0; 
			9'd386:  coeff = 10'sd0; 
			9'd387:  coeff = 10'sd0; 
			9'd388:  coeff = 10'sd0; 
			9'd389:  coeff = 10'sd0; 
			9'd390:  coeff = 10'sd0; 
			9'd391:  coeff = 10'sd0; 
			9'd392:  coeff = 10'sd0; 
			9'd393:  coeff = 10'sd0; 
			9'd394:  coeff = 10'sd0; 
			9'd395:  coeff = 10'sd0; 
			9'd396:  coeff = 10'sd0; 
			9'd397:  coeff = 10'sd0; 
			9'd398:  coeff = 10'sd0; 
			9'd399:  coeff = 10'sd0; 
			9'd400:  coeff = 10'sd0; 

			default: coeff = 10'hXXX;
		endcase
endmodule


module coeffs400tap_600_1200Hz(
  input wire [8:0] index,
  output reg signed [9:0] coeff
);
  // tools will turn this into a 401x10 ROM
	always @(index)
		case (index)
		
			9'd0:  coeff = 10'sd0; 
			9'd1:  coeff = 10'sd0; 
			9'd2:  coeff = 10'sd0; 
			9'd3:  coeff = 10'sd0; 
			9'd4:  coeff = 10'sd0; 
			9'd5:  coeff = 10'sd0; 
			9'd6:  coeff = 10'sd0; 
			9'd7:  coeff = 10'sd0; 
			9'd8:  coeff = 10'sd0; 
			9'd9:  coeff = 10'sd0; 
			9'd10:  coeff = 10'sd0; 
			9'd11:  coeff = 10'sd0; 
			9'd12:  coeff = 10'sd0; 
			9'd13:  coeff = 10'sd0; 
			9'd14:  coeff = 10'sd0; 
			9'd15:  coeff = 10'sd0; 
			9'd16:  coeff = 10'sd0; 
			9'd17:  coeff = 10'sd0; 
			9'd18:  coeff = 10'sd0; 
			9'd19:  coeff = 10'sd0; 
			9'd20:  coeff = 10'sd0; 
			9'd21:  coeff = 10'sd0; 
			9'd22:  coeff = 10'sd0; 
			9'd23:  coeff = 10'sd0; 
			9'd24:  coeff = 10'sd0; 
			9'd25:  coeff = 10'sd0; 
			9'd26:  coeff = 10'sd0; 
			9'd27:  coeff = 10'sd0; 
			9'd28:  coeff = 10'sd0; 
			9'd29:  coeff = 10'sd0; 
			9'd30:  coeff = 10'sd0; 
			9'd31:  coeff = 10'sd0; 
			9'd32:  coeff = 10'sd0; 
			9'd33:  coeff = 10'sd0; 
			9'd34:  coeff = 10'sd0; 
			9'd35:  coeff = 10'sd0; 
			9'd36:  coeff = 10'sd0; 
			9'd37:  coeff = 10'sd0; 
			9'd38:  coeff = 10'sd0; 
			9'd39:  coeff = 10'sd0; 
			9'd40:  coeff = 10'sd0; 
			9'd41:  coeff = 10'sd0; 
			9'd42:  coeff = 10'sd0; 
			9'd43:  coeff = 10'sd0; 
			9'd44:  coeff = 10'sd0; 
			9'd45:  coeff = 10'sd0; 
			9'd46:  coeff = 10'sd0; 
			9'd47:  coeff = 10'sd0; 
			9'd48:  coeff = 10'sd0; 
			9'd49:  coeff = 10'sd0; 
			9'd50:  coeff = 10'sd0; 
			9'd51:  coeff = 10'sd0; 
			9'd52:  coeff = 10'sd0; 
			9'd53:  coeff = 10'sd0; 
			9'd54:  coeff = 10'sd0; 
			9'd55:  coeff = 10'sd0; 
			9'd56:  coeff = 10'sd0; 
			9'd57:  coeff = 10'sd0; 
			9'd58:  coeff = 10'sd0; 
			9'd59:  coeff = 10'sd0; 
			9'd60:  coeff = 10'sd0; 
			9'd61:  coeff = 10'sd0; 
			9'd62:  coeff = 10'sd0; 
			9'd63:  coeff = 10'sd0; 
			9'd64:  coeff = 10'sd0; 
			9'd65:  coeff = 10'sd0; 
			9'd66:  coeff = 10'sd0; 
			9'd67:  coeff = 10'sd0; 
			9'd68:  coeff = 10'sd0; 
			9'd69:  coeff = 10'sd0; 
			9'd70:  coeff = 10'sd0; 
			9'd71:  coeff = 10'sd0; 
			9'd72:  coeff = 10'sd0; 
			9'd73:  coeff = 10'sd0; 
			9'd74:  coeff = 10'sd0; 
			9'd75:  coeff = 10'sd0; 
			9'd76:  coeff = 10'sd0; 
			9'd77:  coeff = 10'sd0; 
			9'd78:  coeff = 10'sd0; 
			9'd79:  coeff = 10'sd0; 
			9'd80:  coeff = 10'sd0; 
			9'd81:  coeff = 10'sd0; 
			9'd82:  coeff = 10'sd0; 
			9'd83:  coeff = 10'sd0; 
			9'd84:  coeff = 10'sd0; 
			9'd85:  coeff = 10'sd0; 
			9'd86:  coeff = -10'sd1; 
			9'd87:  coeff = -10'sd1; 
			9'd88:  coeff = -10'sd1; 
			9'd89:  coeff = -10'sd1; 
			9'd90:  coeff = -10'sd1; 
			9'd91:  coeff = -10'sd1; 
			9'd92:  coeff = -10'sd1; 
			9'd93:  coeff = -10'sd1; 
			9'd94:  coeff = -10'sd1; 
			9'd95:  coeff = -10'sd1; 
			9'd96:  coeff = -10'sd1; 
			9'd97:  coeff = -10'sd1; 
			9'd98:  coeff = -10'sd1; 
			9'd99:  coeff = -10'sd1; 
			9'd100:  coeff = -10'sd1; 
			9'd101:  coeff = -10'sd1; 
			9'd102:  coeff = -10'sd1; 
			9'd103:  coeff = 10'sd0; 
			9'd104:  coeff = 10'sd0; 
			9'd105:  coeff = 10'sd0; 
			9'd106:  coeff = 10'sd0; 
			9'd107:  coeff = 10'sd0; 
			9'd108:  coeff = 10'sd0; 
			9'd109:  coeff = 10'sd0; 
			9'd110:  coeff = 10'sd0; 
			9'd111:  coeff = 10'sd0; 
			9'd112:  coeff = 10'sd0; 
			9'd113:  coeff = 10'sd0; 
			9'd114:  coeff = 10'sd0; 
			9'd115:  coeff = 10'sd0; 
			9'd116:  coeff = 10'sd0; 
			9'd117:  coeff = 10'sd0; 
			9'd118:  coeff = 10'sd0; 
			9'd119:  coeff = 10'sd0; 
			9'd120:  coeff = 10'sd0; 
			9'd121:  coeff = 10'sd0; 
			9'd122:  coeff = 10'sd0; 
			9'd123:  coeff = 10'sd0; 
			9'd124:  coeff = -10'sd1; 
			9'd125:  coeff = -10'sd1; 
			9'd126:  coeff = -10'sd1; 
			9'd127:  coeff = -10'sd1; 
			9'd128:  coeff = -10'sd1; 
			9'd129:  coeff = -10'sd1; 
			9'd130:  coeff = -10'sd1; 
			9'd131:  coeff = -10'sd1; 
			9'd132:  coeff = 10'sd0; 
			9'd133:  coeff = 10'sd0; 
			9'd134:  coeff = 10'sd0; 
			9'd135:  coeff = 10'sd1; 
			9'd136:  coeff = 10'sd1; 
			9'd137:  coeff = 10'sd2; 
			9'd138:  coeff = 10'sd2; 
			9'd139:  coeff = 10'sd3; 
			9'd140:  coeff = 10'sd3; 
			9'd141:  coeff = 10'sd4; 
			9'd142:  coeff = 10'sd5; 
			9'd143:  coeff = 10'sd5; 
			9'd144:  coeff = 10'sd6; 
			9'd145:  coeff = 10'sd6; 
			9'd146:  coeff = 10'sd7; 
			9'd147:  coeff = 10'sd7; 
			9'd148:  coeff = 10'sd8; 
			9'd149:  coeff = 10'sd8; 
			9'd150:  coeff = 10'sd8; 
			9'd151:  coeff = 10'sd8; 
			9'd152:  coeff = 10'sd8; 
			9'd153:  coeff = 10'sd7; 
			9'd154:  coeff = 10'sd7; 
			9'd155:  coeff = 10'sd6; 
			9'd156:  coeff = 10'sd5; 
			9'd157:  coeff = 10'sd4; 
			9'd158:  coeff = 10'sd3; 
			9'd159:  coeff = 10'sd2; 
			9'd160:  coeff = 10'sd0; 
			9'd161:  coeff = -10'sd2; 
			9'd162:  coeff = -10'sd3; 
			9'd163:  coeff = -10'sd5; 
			9'd164:  coeff = -10'sd7; 
			9'd165:  coeff = -10'sd9; 
			9'd166:  coeff = -10'sd10; 
			9'd167:  coeff = -10'sd12; 
			9'd168:  coeff = -10'sd14; 
			9'd169:  coeff = -10'sd15; 
			9'd170:  coeff = -10'sd17; 
			9'd171:  coeff = -10'sd18; 
			9'd172:  coeff = -10'sd19; 
			9'd173:  coeff = -10'sd19; 
			9'd174:  coeff = -10'sd20; 
			9'd175:  coeff = -10'sd20; 
			9'd176:  coeff = -10'sd20; 
			9'd177:  coeff = -10'sd19; 
			9'd178:  coeff = -10'sd18; 
			9'd179:  coeff = -10'sd17; 
			9'd180:  coeff = -10'sd16; 
			9'd181:  coeff = -10'sd14; 
			9'd182:  coeff = -10'sd12; 
			9'd183:  coeff = -10'sd10; 
			9'd184:  coeff = -10'sd7; 
			9'd185:  coeff = -10'sd5; 
			9'd186:  coeff = -10'sd2; 
			9'd187:  coeff = 10'sd1; 
			9'd188:  coeff = 10'sd4; 
			9'd189:  coeff = 10'sd7; 
			9'd190:  coeff = 10'sd10; 
			9'd191:  coeff = 10'sd12; 
			9'd192:  coeff = 10'sd15; 
			9'd193:  coeff = 10'sd17; 
			9'd194:  coeff = 10'sd19; 
			9'd195:  coeff = 10'sd21; 
			9'd196:  coeff = 10'sd23; 
			9'd197:  coeff = 10'sd24; 
			9'd198:  coeff = 10'sd25; 
			9'd199:  coeff = 10'sd26; 
			9'd200:  coeff = 10'sd26; 
			9'd201:  coeff = 10'sd26; 
			9'd202:  coeff = 10'sd25; 
			9'd203:  coeff = 10'sd24; 
			9'd204:  coeff = 10'sd23; 
			9'd205:  coeff = 10'sd21; 
			9'd206:  coeff = 10'sd19; 
			9'd207:  coeff = 10'sd17; 
			9'd208:  coeff = 10'sd15; 
			9'd209:  coeff = 10'sd12; 
			9'd210:  coeff = 10'sd10; 
			9'd211:  coeff = 10'sd7; 
			9'd212:  coeff = 10'sd4; 
			9'd213:  coeff = 10'sd1; 
			9'd214:  coeff = -10'sd2; 
			9'd215:  coeff = -10'sd5; 
			9'd216:  coeff = -10'sd7; 
			9'd217:  coeff = -10'sd10; 
			9'd218:  coeff = -10'sd12; 
			9'd219:  coeff = -10'sd14; 
			9'd220:  coeff = -10'sd16; 
			9'd221:  coeff = -10'sd17; 
			9'd222:  coeff = -10'sd18; 
			9'd223:  coeff = -10'sd19; 
			9'd224:  coeff = -10'sd20; 
			9'd225:  coeff = -10'sd20; 
			9'd226:  coeff = -10'sd20; 
			9'd227:  coeff = -10'sd19; 
			9'd228:  coeff = -10'sd19; 
			9'd229:  coeff = -10'sd18; 
			9'd230:  coeff = -10'sd17; 
			9'd231:  coeff = -10'sd15; 
			9'd232:  coeff = -10'sd14; 
			9'd233:  coeff = -10'sd12; 
			9'd234:  coeff = -10'sd10; 
			9'd235:  coeff = -10'sd9; 
			9'd236:  coeff = -10'sd7; 
			9'd237:  coeff = -10'sd5; 
			9'd238:  coeff = -10'sd3; 
			9'd239:  coeff = -10'sd2; 
			9'd240:  coeff = 10'sd0; 
			9'd241:  coeff = 10'sd2; 
			9'd242:  coeff = 10'sd3; 
			9'd243:  coeff = 10'sd4; 
			9'd244:  coeff = 10'sd5; 
			9'd245:  coeff = 10'sd6; 
			9'd246:  coeff = 10'sd7; 
			9'd247:  coeff = 10'sd7; 
			9'd248:  coeff = 10'sd8; 
			9'd249:  coeff = 10'sd8; 
			9'd250:  coeff = 10'sd8; 
			9'd251:  coeff = 10'sd8; 
			9'd252:  coeff = 10'sd8; 
			9'd253:  coeff = 10'sd7; 
			9'd254:  coeff = 10'sd7; 
			9'd255:  coeff = 10'sd6; 
			9'd256:  coeff = 10'sd6; 
			9'd257:  coeff = 10'sd5; 
			9'd258:  coeff = 10'sd5; 
			9'd259:  coeff = 10'sd4; 
			9'd260:  coeff = 10'sd3; 
			9'd261:  coeff = 10'sd3; 
			9'd262:  coeff = 10'sd2; 
			9'd263:  coeff = 10'sd2; 
			9'd264:  coeff = 10'sd1; 
			9'd265:  coeff = 10'sd1; 
			9'd266:  coeff = 10'sd0; 
			9'd267:  coeff = 10'sd0; 
			9'd268:  coeff = 10'sd0; 
			9'd269:  coeff = -10'sd1; 
			9'd270:  coeff = -10'sd1; 
			9'd271:  coeff = -10'sd1; 
			9'd272:  coeff = -10'sd1; 
			9'd273:  coeff = -10'sd1; 
			9'd274:  coeff = -10'sd1; 
			9'd275:  coeff = -10'sd1; 
			9'd276:  coeff = -10'sd1; 
			9'd277:  coeff = 10'sd0; 
			9'd278:  coeff = 10'sd0; 
			9'd279:  coeff = 10'sd0; 
			9'd280:  coeff = 10'sd0; 
			9'd281:  coeff = 10'sd0; 
			9'd282:  coeff = 10'sd0; 
			9'd283:  coeff = 10'sd0; 
			9'd284:  coeff = 10'sd0; 
			9'd285:  coeff = 10'sd0; 
			9'd286:  coeff = 10'sd0; 
			9'd287:  coeff = 10'sd0; 
			9'd288:  coeff = 10'sd0; 
			9'd289:  coeff = 10'sd0; 
			9'd290:  coeff = 10'sd0; 
			9'd291:  coeff = 10'sd0; 
			9'd292:  coeff = 10'sd0; 
			9'd293:  coeff = 10'sd0; 
			9'd294:  coeff = 10'sd0; 
			9'd295:  coeff = 10'sd0; 
			9'd296:  coeff = 10'sd0; 
			9'd297:  coeff = 10'sd0; 
			9'd298:  coeff = -10'sd1; 
			9'd299:  coeff = -10'sd1; 
			9'd300:  coeff = -10'sd1; 
			9'd301:  coeff = -10'sd1; 
			9'd302:  coeff = -10'sd1; 
			9'd303:  coeff = -10'sd1; 
			9'd304:  coeff = -10'sd1; 
			9'd305:  coeff = -10'sd1; 
			9'd306:  coeff = -10'sd1; 
			9'd307:  coeff = -10'sd1; 
			9'd308:  coeff = -10'sd1; 
			9'd309:  coeff = -10'sd1; 
			9'd310:  coeff = -10'sd1; 
			9'd311:  coeff = -10'sd1; 
			9'd312:  coeff = -10'sd1; 
			9'd313:  coeff = -10'sd1; 
			9'd314:  coeff = -10'sd1; 
			9'd315:  coeff = 10'sd0; 
			9'd316:  coeff = 10'sd0; 
			9'd317:  coeff = 10'sd0; 
			9'd318:  coeff = 10'sd0; 
			9'd319:  coeff = 10'sd0; 
			9'd320:  coeff = 10'sd0; 
			9'd321:  coeff = 10'sd0; 
			9'd322:  coeff = 10'sd0; 
			9'd323:  coeff = 10'sd0; 
			9'd324:  coeff = 10'sd0; 
			9'd325:  coeff = 10'sd0; 
			9'd326:  coeff = 10'sd0; 
			9'd327:  coeff = 10'sd0; 
			9'd328:  coeff = 10'sd0; 
			9'd329:  coeff = 10'sd0; 
			9'd330:  coeff = 10'sd0; 
			9'd331:  coeff = 10'sd0; 
			9'd332:  coeff = 10'sd0; 
			9'd333:  coeff = 10'sd0; 
			9'd334:  coeff = 10'sd0; 
			9'd335:  coeff = 10'sd0; 
			9'd336:  coeff = 10'sd0; 
			9'd337:  coeff = 10'sd0; 
			9'd338:  coeff = 10'sd0; 
			9'd339:  coeff = 10'sd0; 
			9'd340:  coeff = 10'sd0; 
			9'd341:  coeff = 10'sd0; 
			9'd342:  coeff = 10'sd0; 
			9'd343:  coeff = 10'sd0; 
			9'd344:  coeff = 10'sd0; 
			9'd345:  coeff = 10'sd0; 
			9'd346:  coeff = 10'sd0; 
			9'd347:  coeff = 10'sd0; 
			9'd348:  coeff = 10'sd0; 
			9'd349:  coeff = 10'sd0; 
			9'd350:  coeff = 10'sd0; 
			9'd351:  coeff = 10'sd0; 
			9'd352:  coeff = 10'sd0; 
			9'd353:  coeff = 10'sd0; 
			9'd354:  coeff = 10'sd0; 
			9'd355:  coeff = 10'sd0; 
			9'd356:  coeff = 10'sd0; 
			9'd357:  coeff = 10'sd0; 
			9'd358:  coeff = 10'sd0; 
			9'd359:  coeff = 10'sd0; 
			9'd360:  coeff = 10'sd0; 
			9'd361:  coeff = 10'sd0; 
			9'd362:  coeff = 10'sd0; 
			9'd363:  coeff = 10'sd0; 
			9'd364:  coeff = 10'sd0; 
			9'd365:  coeff = 10'sd0; 
			9'd366:  coeff = 10'sd0; 
			9'd367:  coeff = 10'sd0; 
			9'd368:  coeff = 10'sd0; 
			9'd369:  coeff = 10'sd0; 
			9'd370:  coeff = 10'sd0; 
			9'd371:  coeff = 10'sd0; 
			9'd372:  coeff = 10'sd0; 
			9'd373:  coeff = 10'sd0; 
			9'd374:  coeff = 10'sd0; 
			9'd375:  coeff = 10'sd0; 
			9'd376:  coeff = 10'sd0; 
			9'd377:  coeff = 10'sd0; 
			9'd378:  coeff = 10'sd0; 
			9'd379:  coeff = 10'sd0; 
			9'd380:  coeff = 10'sd0; 
			9'd381:  coeff = 10'sd0; 
			9'd382:  coeff = 10'sd0; 
			9'd383:  coeff = 10'sd0; 
			9'd384:  coeff = 10'sd0; 
			9'd385:  coeff = 10'sd0; 
			9'd386:  coeff = 10'sd0; 
			9'd387:  coeff = 10'sd0; 
			9'd388:  coeff = 10'sd0; 
			9'd389:  coeff = 10'sd0; 
			9'd390:  coeff = 10'sd0; 
			9'd391:  coeff = 10'sd0; 
			9'd392:  coeff = 10'sd0; 
			9'd393:  coeff = 10'sd0; 
			9'd394:  coeff = 10'sd0; 
			9'd395:  coeff = 10'sd0; 
			9'd396:  coeff = 10'sd0; 
			9'd397:  coeff = 10'sd0; 
			9'd398:  coeff = 10'sd0; 
			9'd399:  coeff = 10'sd0; 
			9'd400:  coeff = 10'sd0; 

			default: coeff = 10'hXXX;
		endcase
endmodule


module coeffs400tap_1200_4kHz(
  input wire [8:0] index,
  output reg signed [9:0] coeff
);
  // tools will turn this into a 400x10 ROM
	always @(index)
		case (index)

			9'd0:  coeff = 10'sd0; 
			9'd1:  coeff = 10'sd0; 
			9'd2:  coeff = 10'sd0; 
			9'd3:  coeff = 10'sd0; 
			9'd4:  coeff = 10'sd0; 
			9'd5:  coeff = 10'sd0; 
			9'd6:  coeff = 10'sd0; 
			9'd7:  coeff = 10'sd0; 
			9'd8:  coeff = 10'sd0; 
			9'd9:  coeff = 10'sd0; 
			9'd10:  coeff = 10'sd0; 
			9'd11:  coeff = 10'sd0; 
			9'd12:  coeff = 10'sd0; 
			9'd13:  coeff = 10'sd0; 
			9'd14:  coeff = 10'sd0; 
			9'd15:  coeff = 10'sd0; 
			9'd16:  coeff = 10'sd0; 
			9'd17:  coeff = 10'sd0; 
			9'd18:  coeff = 10'sd0; 
			9'd19:  coeff = 10'sd0; 
			9'd20:  coeff = 10'sd0; 
			9'd21:  coeff = 10'sd0; 
			9'd22:  coeff = 10'sd0; 
			9'd23:  coeff = 10'sd0; 
			9'd24:  coeff = 10'sd0; 
			9'd25:  coeff = 10'sd0; 
			9'd26:  coeff = 10'sd0; 
			9'd27:  coeff = 10'sd0; 
			9'd28:  coeff = 10'sd0; 
			9'd29:  coeff = 10'sd0; 
			9'd30:  coeff = 10'sd0; 
			9'd31:  coeff = 10'sd0; 
			9'd32:  coeff = 10'sd0; 
			9'd33:  coeff = 10'sd0; 
			9'd34:  coeff = 10'sd0; 
			9'd35:  coeff = 10'sd0; 
			9'd36:  coeff = 10'sd0; 
			9'd37:  coeff = 10'sd0; 
			9'd38:  coeff = 10'sd0; 
			9'd39:  coeff = 10'sd0; 
			9'd40:  coeff = 10'sd0; 
			9'd41:  coeff = 10'sd0; 
			9'd42:  coeff = 10'sd0; 
			9'd43:  coeff = 10'sd0; 
			9'd44:  coeff = 10'sd0; 
			9'd45:  coeff = 10'sd0; 
			9'd46:  coeff = 10'sd0; 
			9'd47:  coeff = 10'sd0; 
			9'd48:  coeff = 10'sd0; 
			9'd49:  coeff = 10'sd0; 
			9'd50:  coeff = 10'sd0; 
			9'd51:  coeff = 10'sd0; 
			9'd52:  coeff = 10'sd0; 
			9'd53:  coeff = 10'sd0; 
			9'd54:  coeff = 10'sd0; 
			9'd55:  coeff = 10'sd0; 
			9'd56:  coeff = 10'sd0; 
			9'd57:  coeff = 10'sd0; 
			9'd58:  coeff = 10'sd0; 
			9'd59:  coeff = 10'sd0; 
			9'd60:  coeff = 10'sd0; 
			9'd61:  coeff = 10'sd0; 
			9'd62:  coeff = 10'sd0; 
			9'd63:  coeff = 10'sd0; 
			9'd64:  coeff = 10'sd0; 
			9'd65:  coeff = 10'sd0; 
			9'd66:  coeff = 10'sd0; 
			9'd67:  coeff = 10'sd0; 
			9'd68:  coeff = 10'sd0; 
			9'd69:  coeff = 10'sd0; 
			9'd70:  coeff = 10'sd0; 
			9'd71:  coeff = 10'sd0; 
			9'd72:  coeff = 10'sd0; 
			9'd73:  coeff = 10'sd0; 
			9'd74:  coeff = 10'sd0; 
			9'd75:  coeff = 10'sd0; 
			9'd76:  coeff = 10'sd0; 
			9'd77:  coeff = 10'sd0; 
			9'd78:  coeff = 10'sd0; 
			9'd79:  coeff = 10'sd0; 
			9'd80:  coeff = 10'sd0; 
			9'd81:  coeff = 10'sd0; 
			9'd82:  coeff = 10'sd0; 
			9'd83:  coeff = 10'sd0; 
			9'd84:  coeff = 10'sd0; 
			9'd85:  coeff = 10'sd0; 
			9'd86:  coeff = 10'sd0; 
			9'd87:  coeff = 10'sd0; 
			9'd88:  coeff = 10'sd0; 
			9'd89:  coeff = 10'sd0; 
			9'd90:  coeff = 10'sd0; 
			9'd91:  coeff = -10'sd1; 
			9'd92:  coeff = -10'sd1; 
			9'd93:  coeff = 10'sd0; 
			9'd94:  coeff = 10'sd0; 
			9'd95:  coeff = 10'sd0; 
			9'd96:  coeff = 10'sd1; 
			9'd97:  coeff = 10'sd1; 
			9'd98:  coeff = 10'sd1; 
			9'd99:  coeff = 10'sd0; 
			9'd100:  coeff = 10'sd0; 
			9'd101:  coeff = 10'sd0; 
			9'd102:  coeff = -10'sd1; 
			9'd103:  coeff = -10'sd1; 
			9'd104:  coeff = -10'sd1; 
			9'd105:  coeff = 10'sd0; 
			9'd106:  coeff = 10'sd0; 
			9'd107:  coeff = 10'sd1; 
			9'd108:  coeff = 10'sd1; 
			9'd109:  coeff = 10'sd1; 
			9'd110:  coeff = 10'sd1; 
			9'd111:  coeff = 10'sd0; 
			9'd112:  coeff = 10'sd0; 
			9'd113:  coeff = -10'sd1; 
			9'd114:  coeff = -10'sd1; 
			9'd115:  coeff = -10'sd1; 
			9'd116:  coeff = -10'sd1; 
			9'd117:  coeff = -10'sd1; 
			9'd118:  coeff = 10'sd0; 
			9'd119:  coeff = 10'sd1; 
			9'd120:  coeff = 10'sd2; 
			9'd121:  coeff = 10'sd2; 
			9'd122:  coeff = 10'sd1; 
			9'd123:  coeff = 10'sd1; 
			9'd124:  coeff = 10'sd0; 
			9'd125:  coeff = -10'sd1; 
			9'd126:  coeff = -10'sd2; 
			9'd127:  coeff = -10'sd2; 
			9'd128:  coeff = -10'sd2; 
			9'd129:  coeff = 10'sd0; 
			9'd130:  coeff = 10'sd1; 
			9'd131:  coeff = 10'sd2; 
			9'd132:  coeff = 10'sd2; 
			9'd133:  coeff = 10'sd2; 
			9'd134:  coeff = 10'sd2; 
			9'd135:  coeff = 10'sd0; 
			9'd136:  coeff = -10'sd1; 
			9'd137:  coeff = -10'sd2; 
			9'd138:  coeff = -10'sd3; 
			9'd139:  coeff = -10'sd3; 
			9'd140:  coeff = -10'sd2; 
			9'd141:  coeff = 10'sd0; 
			9'd142:  coeff = 10'sd2; 
			9'd143:  coeff = 10'sd3; 
			9'd144:  coeff = 10'sd4; 
			9'd145:  coeff = 10'sd3; 
			9'd146:  coeff = 10'sd2; 
			9'd147:  coeff = 10'sd0; 
			9'd148:  coeff = -10'sd2; 
			9'd149:  coeff = -10'sd4; 
			9'd150:  coeff = -10'sd5; 
			9'd151:  coeff = -10'sd4; 
			9'd152:  coeff = -10'sd2; 
			9'd153:  coeff = 10'sd0; 
			9'd154:  coeff = 10'sd3; 
			9'd155:  coeff = 10'sd5; 
			9'd156:  coeff = 10'sd6; 
			9'd157:  coeff = 10'sd5; 
			9'd158:  coeff = 10'sd3; 
			9'd159:  coeff = -10'sd1; 
			9'd160:  coeff = -10'sd4; 
			9'd161:  coeff = -10'sd6; 
			9'd162:  coeff = -10'sd7; 
			9'd163:  coeff = -10'sd6; 
			9'd164:  coeff = -10'sd3; 
			9'd165:  coeff = 10'sd1; 
			9'd166:  coeff = 10'sd5; 
			9'd167:  coeff = 10'sd8; 
			9'd168:  coeff = 10'sd9; 
			9'd169:  coeff = 10'sd7; 
			9'd170:  coeff = 10'sd3; 
			9'd171:  coeff = -10'sd2; 
			9'd172:  coeff = -10'sd7; 
			9'd173:  coeff = -10'sd11; 
			9'd174:  coeff = -10'sd11; 
			9'd175:  coeff = -10'sd8; 
			9'd176:  coeff = -10'sd3; 
			9'd177:  coeff = 10'sd4; 
			9'd178:  coeff = 10'sd10; 
			9'd179:  coeff = 10'sd14; 
			9'd180:  coeff = 10'sd15; 
			9'd181:  coeff = 10'sd11; 
			9'd182:  coeff = 10'sd3; 
			9'd183:  coeff = -10'sd6; 
			9'd184:  coeff = -10'sd15; 
			9'd185:  coeff = -10'sd21; 
			9'd186:  coeff = -10'sd21; 
			9'd187:  coeff = -10'sd15; 
			9'd188:  coeff = -10'sd3; 
			9'd189:  coeff = 10'sd12; 
			9'd190:  coeff = 10'sd26; 
			9'd191:  coeff = 10'sd36; 
			9'd192:  coeff = 10'sd37; 
			9'd193:  coeff = 10'sd26; 
			9'd194:  coeff = 10'sd3; 
			9'd195:  coeff = -10'sd29; 
			9'd196:  coeff = -10'sd69; 
			9'd197:  coeff = -10'sd108; 
			9'd198:  coeff = -10'sd143; 
			9'd199:  coeff = -10'sd166; 
			9'd200:  coeff = 10'sd850; 
			9'd201:  coeff = -10'sd166; 
			9'd202:  coeff = -10'sd143; 
			9'd203:  coeff = -10'sd108; 
			9'd204:  coeff = -10'sd69; 
			9'd205:  coeff = -10'sd29; 
			9'd206:  coeff = 10'sd3; 
			9'd207:  coeff = 10'sd26; 
			9'd208:  coeff = 10'sd37; 
			9'd209:  coeff = 10'sd36; 
			9'd210:  coeff = 10'sd26; 
			9'd211:  coeff = 10'sd12; 
			9'd212:  coeff = -10'sd3; 
			9'd213:  coeff = -10'sd15; 
			9'd214:  coeff = -10'sd21; 
			9'd215:  coeff = -10'sd21; 
			9'd216:  coeff = -10'sd15; 
			9'd217:  coeff = -10'sd6; 
			9'd218:  coeff = 10'sd3; 
			9'd219:  coeff = 10'sd11; 
			9'd220:  coeff = 10'sd15; 
			9'd221:  coeff = 10'sd14; 
			9'd222:  coeff = 10'sd10; 
			9'd223:  coeff = 10'sd4; 
			9'd224:  coeff = -10'sd3; 
			9'd225:  coeff = -10'sd8; 
			9'd226:  coeff = -10'sd11; 
			9'd227:  coeff = -10'sd11; 
			9'd228:  coeff = -10'sd7; 
			9'd229:  coeff = -10'sd2; 
			9'd230:  coeff = 10'sd3; 
			9'd231:  coeff = 10'sd7; 
			9'd232:  coeff = 10'sd9; 
			9'd233:  coeff = 10'sd8; 
			9'd234:  coeff = 10'sd5; 
			9'd235:  coeff = 10'sd1; 
			9'd236:  coeff = -10'sd3; 
			9'd237:  coeff = -10'sd6; 
			9'd238:  coeff = -10'sd7; 
			9'd239:  coeff = -10'sd6; 
			9'd240:  coeff = -10'sd4; 
			9'd241:  coeff = -10'sd1; 
			9'd242:  coeff = 10'sd3; 
			9'd243:  coeff = 10'sd5; 
			9'd244:  coeff = 10'sd6; 
			9'd245:  coeff = 10'sd5; 
			9'd246:  coeff = 10'sd3; 
			9'd247:  coeff = 10'sd0; 
			9'd248:  coeff = -10'sd2; 
			9'd249:  coeff = -10'sd4; 
			9'd250:  coeff = -10'sd5; 
			9'd251:  coeff = -10'sd4; 
			9'd252:  coeff = -10'sd2; 
			9'd253:  coeff = 10'sd0; 
			9'd254:  coeff = 10'sd2; 
			9'd255:  coeff = 10'sd3; 
			9'd256:  coeff = 10'sd4; 
			9'd257:  coeff = 10'sd3; 
			9'd258:  coeff = 10'sd2; 
			9'd259:  coeff = 10'sd0; 
			9'd260:  coeff = -10'sd2; 
			9'd261:  coeff = -10'sd3; 
			9'd262:  coeff = -10'sd3; 
			9'd263:  coeff = -10'sd2; 
			9'd264:  coeff = -10'sd1; 
			9'd265:  coeff = 10'sd0; 
			9'd266:  coeff = 10'sd2; 
			9'd267:  coeff = 10'sd2; 
			9'd268:  coeff = 10'sd2; 
			9'd269:  coeff = 10'sd2; 
			9'd270:  coeff = 10'sd1; 
			9'd271:  coeff = 10'sd0; 
			9'd272:  coeff = -10'sd2; 
			9'd273:  coeff = -10'sd2; 
			9'd274:  coeff = -10'sd2; 
			9'd275:  coeff = -10'sd1; 
			9'd276:  coeff = 10'sd0; 
			9'd277:  coeff = 10'sd1; 
			9'd278:  coeff = 10'sd1; 
			9'd279:  coeff = 10'sd2; 
			9'd280:  coeff = 10'sd2; 
			9'd281:  coeff = 10'sd1; 
			9'd282:  coeff = 10'sd0; 
			9'd283:  coeff = -10'sd1; 
			9'd284:  coeff = -10'sd1; 
			9'd285:  coeff = -10'sd1; 
			9'd286:  coeff = -10'sd1; 
			9'd287:  coeff = -10'sd1; 
			9'd288:  coeff = 10'sd0; 
			9'd289:  coeff = 10'sd0; 
			9'd290:  coeff = 10'sd1; 
			9'd291:  coeff = 10'sd1; 
			9'd292:  coeff = 10'sd1; 
			9'd293:  coeff = 10'sd1; 
			9'd294:  coeff = 10'sd0; 
			9'd295:  coeff = 10'sd0; 
			9'd296:  coeff = -10'sd1; 
			9'd297:  coeff = -10'sd1; 
			9'd298:  coeff = -10'sd1; 
			9'd299:  coeff = 10'sd0; 
			9'd300:  coeff = 10'sd0; 
			9'd301:  coeff = 10'sd0; 
			9'd302:  coeff = 10'sd1; 
			9'd303:  coeff = 10'sd1; 
			9'd304:  coeff = 10'sd1; 
			9'd305:  coeff = 10'sd0; 
			9'd306:  coeff = 10'sd0; 
			9'd307:  coeff = 10'sd0; 
			9'd308:  coeff = -10'sd1; 
			9'd309:  coeff = -10'sd1; 
			9'd310:  coeff = 10'sd0; 
			9'd311:  coeff = 10'sd0; 
			9'd312:  coeff = 10'sd0; 
			9'd313:  coeff = 10'sd0; 
			9'd314:  coeff = 10'sd0; 
			9'd315:  coeff = 10'sd0; 
			9'd316:  coeff = 10'sd0; 
			9'd317:  coeff = 10'sd0; 
			9'd318:  coeff = 10'sd0; 
			9'd319:  coeff = 10'sd0; 
			9'd320:  coeff = 10'sd0; 
			9'd321:  coeff = 10'sd0; 
			9'd322:  coeff = 10'sd0; 
			9'd323:  coeff = 10'sd0; 
			9'd324:  coeff = 10'sd0; 
			9'd325:  coeff = 10'sd0; 
			9'd326:  coeff = 10'sd0; 
			9'd327:  coeff = 10'sd0; 
			9'd328:  coeff = 10'sd0; 
			9'd329:  coeff = 10'sd0; 
			9'd330:  coeff = 10'sd0; 
			9'd331:  coeff = 10'sd0; 
			9'd332:  coeff = 10'sd0; 
			9'd333:  coeff = 10'sd0; 
			9'd334:  coeff = 10'sd0; 
			9'd335:  coeff = 10'sd0; 
			9'd336:  coeff = 10'sd0; 
			9'd337:  coeff = 10'sd0; 
			9'd338:  coeff = 10'sd0; 
			9'd339:  coeff = 10'sd0; 
			9'd340:  coeff = 10'sd0; 
			9'd341:  coeff = 10'sd0; 
			9'd342:  coeff = 10'sd0; 
			9'd343:  coeff = 10'sd0; 
			9'd344:  coeff = 10'sd0; 
			9'd345:  coeff = 10'sd0; 
			9'd346:  coeff = 10'sd0; 
			9'd347:  coeff = 10'sd0; 
			9'd348:  coeff = 10'sd0; 
			9'd349:  coeff = 10'sd0; 
			9'd350:  coeff = 10'sd0; 
			9'd351:  coeff = 10'sd0; 
			9'd352:  coeff = 10'sd0; 
			9'd353:  coeff = 10'sd0; 
			9'd354:  coeff = 10'sd0; 
			9'd355:  coeff = 10'sd0; 
			9'd356:  coeff = 10'sd0; 
			9'd357:  coeff = 10'sd0; 
			9'd358:  coeff = 10'sd0; 
			9'd359:  coeff = 10'sd0; 
			9'd360:  coeff = 10'sd0; 
			9'd361:  coeff = 10'sd0; 
			9'd362:  coeff = 10'sd0; 
			9'd363:  coeff = 10'sd0; 
			9'd364:  coeff = 10'sd0; 
			9'd365:  coeff = 10'sd0; 
			9'd366:  coeff = 10'sd0; 
			9'd367:  coeff = 10'sd0; 
			9'd368:  coeff = 10'sd0; 
			9'd369:  coeff = 10'sd0; 
			9'd370:  coeff = 10'sd0; 
			9'd371:  coeff = 10'sd0; 
			9'd372:  coeff = 10'sd0; 
			9'd373:  coeff = 10'sd0; 
			9'd374:  coeff = 10'sd0; 
			9'd375:  coeff = 10'sd0; 
			9'd376:  coeff = 10'sd0; 
			9'd377:  coeff = 10'sd0; 
			9'd378:  coeff = 10'sd0; 
			9'd379:  coeff = 10'sd0; 
			9'd380:  coeff = 10'sd0; 
			9'd381:  coeff = 10'sd0; 
			9'd382:  coeff = 10'sd0; 
			9'd383:  coeff = 10'sd0; 
			9'd384:  coeff = 10'sd0; 
			9'd385:  coeff = 10'sd0; 
			9'd386:  coeff = 10'sd0; 
			9'd387:  coeff = 10'sd0; 
			9'd388:  coeff = 10'sd0; 
			9'd389:  coeff = 10'sd0; 
			9'd390:  coeff = 10'sd0; 
			9'd391:  coeff = 10'sd0; 
			9'd392:  coeff = 10'sd0; 
			9'd393:  coeff = 10'sd0; 
			9'd394:  coeff = 10'sd0; 
			9'd395:  coeff = 10'sd0; 
			9'd396:  coeff = 10'sd0; 
			9'd397:  coeff = 10'sd0; 
			9'd398:  coeff = 10'sd0; 
			9'd399:  coeff = 10'sd0; 
			9'd400:  coeff = 10'sd0; 

			default: coeff = 10'hXXX;
		endcase
endmodule


module coeffs400tap_above_4kHz(
  input wire [8:0] index,
  output reg signed [9:0] coeff
);
  // tools will turn this into a 401x10 ROM
	always @(index)
		case (index)

			9'd0:  coeff = 10'sd0; 
			9'd1:  coeff = 10'sd0; 
			9'd2:  coeff = 10'sd0; 
			9'd3:  coeff = 10'sd0; 
			9'd4:  coeff = 10'sd0; 
			9'd5:  coeff = 10'sd0; 
			9'd6:  coeff = 10'sd0; 
			9'd7:  coeff = 10'sd0; 
			9'd8:  coeff = 10'sd0; 
			9'd9:  coeff = 10'sd0; 
			9'd10:  coeff = 10'sd0; 
			9'd11:  coeff = 10'sd0; 
			9'd12:  coeff = 10'sd0; 
			9'd13:  coeff = 10'sd0; 
			9'd14:  coeff = 10'sd0; 
			9'd15:  coeff = 10'sd0; 
			9'd16:  coeff = 10'sd0; 
			9'd17:  coeff = 10'sd0; 
			9'd18:  coeff = 10'sd0; 
			9'd19:  coeff = 10'sd0; 
			9'd20:  coeff = 10'sd0; 
			9'd21:  coeff = 10'sd0; 
			9'd22:  coeff = 10'sd0; 
			9'd23:  coeff = 10'sd0; 
			9'd24:  coeff = 10'sd0; 
			9'd25:  coeff = 10'sd0; 
			9'd26:  coeff = 10'sd0; 
			9'd27:  coeff = 10'sd0; 
			9'd28:  coeff = 10'sd0; 
			9'd29:  coeff = 10'sd0; 
			9'd30:  coeff = 10'sd0; 
			9'd31:  coeff = 10'sd0; 
			9'd32:  coeff = 10'sd0; 
			9'd33:  coeff = 10'sd0; 
			9'd34:  coeff = 10'sd0; 
			9'd35:  coeff = 10'sd0; 
			9'd36:  coeff = 10'sd0; 
			9'd37:  coeff = 10'sd0; 
			9'd38:  coeff = 10'sd0; 
			9'd39:  coeff = 10'sd0; 
			9'd40:  coeff = 10'sd0; 
			9'd41:  coeff = 10'sd0; 
			9'd42:  coeff = 10'sd0; 
			9'd43:  coeff = 10'sd0; 
			9'd44:  coeff = 10'sd0; 
			9'd45:  coeff = 10'sd0; 
			9'd46:  coeff = 10'sd0; 
			9'd47:  coeff = 10'sd0; 
			9'd48:  coeff = 10'sd0; 
			9'd49:  coeff = 10'sd0; 
			9'd50:  coeff = 10'sd0; 
			9'd51:  coeff = 10'sd0; 
			9'd52:  coeff = 10'sd0; 
			9'd53:  coeff = 10'sd0; 
			9'd54:  coeff = 10'sd0; 
			9'd55:  coeff = 10'sd0; 
			9'd56:  coeff = 10'sd0; 
			9'd57:  coeff = 10'sd0; 
			9'd58:  coeff = 10'sd0; 
			9'd59:  coeff = 10'sd0; 
			9'd60:  coeff = 10'sd0; 
			9'd61:  coeff = 10'sd0; 
			9'd62:  coeff = 10'sd0; 
			9'd63:  coeff = 10'sd0; 
			9'd64:  coeff = 10'sd0; 
			9'd65:  coeff = 10'sd0; 
			9'd66:  coeff = 10'sd0; 
			9'd67:  coeff = 10'sd0; 
			9'd68:  coeff = 10'sd0; 
			9'd69:  coeff = 10'sd0; 
			9'd70:  coeff = 10'sd0; 
			9'd71:  coeff = 10'sd0; 
			9'd72:  coeff = 10'sd0; 
			9'd73:  coeff = 10'sd0; 
			9'd74:  coeff = 10'sd0; 
			9'd75:  coeff = 10'sd0; 
			9'd76:  coeff = 10'sd0; 
			9'd77:  coeff = 10'sd0; 
			9'd78:  coeff = 10'sd0; 
			9'd79:  coeff = 10'sd0; 
			9'd80:  coeff = 10'sd0; 
			9'd81:  coeff = 10'sd0; 
			9'd82:  coeff = 10'sd0; 
			9'd83:  coeff = 10'sd0; 
			9'd84:  coeff = 10'sd0; 
			9'd85:  coeff = 10'sd0; 
			9'd86:  coeff = 10'sd0; 
			9'd87:  coeff = 10'sd0; 
			9'd88:  coeff = 10'sd0; 
			9'd89:  coeff = 10'sd0; 
			9'd90:  coeff = 10'sd0; 
			9'd91:  coeff = -10'sd1; 
			9'd92:  coeff = -10'sd1; 
			9'd93:  coeff = 10'sd0; 
			9'd94:  coeff = 10'sd0; 
			9'd95:  coeff = 10'sd0; 
			9'd96:  coeff = 10'sd1; 
			9'd97:  coeff = 10'sd1; 
			9'd98:  coeff = 10'sd1; 
			9'd99:  coeff = 10'sd0; 
			9'd100:  coeff = 10'sd0; 
			9'd101:  coeff = 10'sd0; 
			9'd102:  coeff = -10'sd1; 
			9'd103:  coeff = -10'sd1; 
			9'd104:  coeff = -10'sd1; 
			9'd105:  coeff = 10'sd0; 
			9'd106:  coeff = 10'sd0; 
			9'd107:  coeff = 10'sd1; 
			9'd108:  coeff = 10'sd1; 
			9'd109:  coeff = 10'sd1; 
			9'd110:  coeff = 10'sd1; 
			9'd111:  coeff = 10'sd0; 
			9'd112:  coeff = 10'sd0; 
			9'd113:  coeff = -10'sd1; 
			9'd114:  coeff = -10'sd1; 
			9'd115:  coeff = -10'sd1; 
			9'd116:  coeff = -10'sd1; 
			9'd117:  coeff = -10'sd1; 
			9'd118:  coeff = 10'sd0; 
			9'd119:  coeff = 10'sd1; 
			9'd120:  coeff = 10'sd2; 
			9'd121:  coeff = 10'sd2; 
			9'd122:  coeff = 10'sd1; 
			9'd123:  coeff = 10'sd1; 
			9'd124:  coeff = 10'sd0; 
			9'd125:  coeff = -10'sd1; 
			9'd126:  coeff = -10'sd2; 
			9'd127:  coeff = -10'sd2; 
			9'd128:  coeff = -10'sd2; 
			9'd129:  coeff = 10'sd0; 
			9'd130:  coeff = 10'sd1; 
			9'd131:  coeff = 10'sd2; 
			9'd132:  coeff = 10'sd2; 
			9'd133:  coeff = 10'sd2; 
			9'd134:  coeff = 10'sd2; 
			9'd135:  coeff = 10'sd0; 
			9'd136:  coeff = -10'sd1; 
			9'd137:  coeff = -10'sd2; 
			9'd138:  coeff = -10'sd3; 
			9'd139:  coeff = -10'sd3; 
			9'd140:  coeff = -10'sd2; 
			9'd141:  coeff = 10'sd0; 
			9'd142:  coeff = 10'sd2; 
			9'd143:  coeff = 10'sd3; 
			9'd144:  coeff = 10'sd4; 
			9'd145:  coeff = 10'sd3; 
			9'd146:  coeff = 10'sd2; 
			9'd147:  coeff = 10'sd0; 
			9'd148:  coeff = -10'sd2; 
			9'd149:  coeff = -10'sd4; 
			9'd150:  coeff = -10'sd5; 
			9'd151:  coeff = -10'sd4; 
			9'd152:  coeff = -10'sd2; 
			9'd153:  coeff = 10'sd0; 
			9'd154:  coeff = 10'sd3; 
			9'd155:  coeff = 10'sd5; 
			9'd156:  coeff = 10'sd6; 
			9'd157:  coeff = 10'sd5; 
			9'd158:  coeff = 10'sd3; 
			9'd159:  coeff = -10'sd1; 
			9'd160:  coeff = -10'sd4; 
			9'd161:  coeff = -10'sd6; 
			9'd162:  coeff = -10'sd7; 
			9'd163:  coeff = -10'sd6; 
			9'd164:  coeff = -10'sd3; 
			9'd165:  coeff = 10'sd1; 
			9'd166:  coeff = 10'sd5; 
			9'd167:  coeff = 10'sd8; 
			9'd168:  coeff = 10'sd9; 
			9'd169:  coeff = 10'sd7; 
			9'd170:  coeff = 10'sd3; 
			9'd171:  coeff = -10'sd2; 
			9'd172:  coeff = -10'sd7; 
			9'd173:  coeff = -10'sd11; 
			9'd174:  coeff = -10'sd11; 
			9'd175:  coeff = -10'sd8; 
			9'd176:  coeff = -10'sd3; 
			9'd177:  coeff = 10'sd4; 
			9'd178:  coeff = 10'sd10; 
			9'd179:  coeff = 10'sd14; 
			9'd180:  coeff = 10'sd15; 
			9'd181:  coeff = 10'sd11; 
			9'd182:  coeff = 10'sd3; 
			9'd183:  coeff = -10'sd6; 
			9'd184:  coeff = -10'sd15; 
			9'd185:  coeff = -10'sd21; 
			9'd186:  coeff = -10'sd21; 
			9'd187:  coeff = -10'sd15; 
			9'd188:  coeff = -10'sd3; 
			9'd189:  coeff = 10'sd12; 
			9'd190:  coeff = 10'sd26; 
			9'd191:  coeff = 10'sd36; 
			9'd192:  coeff = 10'sd37; 
			9'd193:  coeff = 10'sd26; 
			9'd194:  coeff = 10'sd3; 
			9'd195:  coeff = -10'sd29; 
			9'd196:  coeff = -10'sd69; 
			9'd197:  coeff = -10'sd108; 
			9'd198:  coeff = -10'sd143; 
			9'd199:  coeff = -10'sd166; 
			9'd200:  coeff = 10'sd850; 
			9'd201:  coeff = -10'sd166; 
			9'd202:  coeff = -10'sd143; 
			9'd203:  coeff = -10'sd108; 
			9'd204:  coeff = -10'sd69; 
			9'd205:  coeff = -10'sd29; 
			9'd206:  coeff = 10'sd3; 
			9'd207:  coeff = 10'sd26; 
			9'd208:  coeff = 10'sd37; 
			9'd209:  coeff = 10'sd36; 
			9'd210:  coeff = 10'sd26; 
			9'd211:  coeff = 10'sd12; 
			9'd212:  coeff = -10'sd3; 
			9'd213:  coeff = -10'sd15; 
			9'd214:  coeff = -10'sd21; 
			9'd215:  coeff = -10'sd21; 
			9'd216:  coeff = -10'sd15; 
			9'd217:  coeff = -10'sd6; 
			9'd218:  coeff = 10'sd3; 
			9'd219:  coeff = 10'sd11; 
			9'd220:  coeff = 10'sd15; 
			9'd221:  coeff = 10'sd14; 
			9'd222:  coeff = 10'sd10; 
			9'd223:  coeff = 10'sd4; 
			9'd224:  coeff = -10'sd3; 
			9'd225:  coeff = -10'sd8; 
			9'd226:  coeff = -10'sd11; 
			9'd227:  coeff = -10'sd11; 
			9'd228:  coeff = -10'sd7; 
			9'd229:  coeff = -10'sd2; 
			9'd230:  coeff = 10'sd3; 
			9'd231:  coeff = 10'sd7; 
			9'd232:  coeff = 10'sd9; 
			9'd233:  coeff = 10'sd8; 
			9'd234:  coeff = 10'sd5; 
			9'd235:  coeff = 10'sd1; 
			9'd236:  coeff = -10'sd3; 
			9'd237:  coeff = -10'sd6; 
			9'd238:  coeff = -10'sd7; 
			9'd239:  coeff = -10'sd6; 
			9'd240:  coeff = -10'sd4; 
			9'd241:  coeff = -10'sd1; 
			9'd242:  coeff = 10'sd3; 
			9'd243:  coeff = 10'sd5; 
			9'd244:  coeff = 10'sd6; 
			9'd245:  coeff = 10'sd5; 
			9'd246:  coeff = 10'sd3; 
			9'd247:  coeff = 10'sd0; 
			9'd248:  coeff = -10'sd2; 
			9'd249:  coeff = -10'sd4; 
			9'd250:  coeff = -10'sd5; 
			9'd251:  coeff = -10'sd4; 
			9'd252:  coeff = -10'sd2; 
			9'd253:  coeff = 10'sd0; 
			9'd254:  coeff = 10'sd2; 
			9'd255:  coeff = 10'sd3; 
			9'd256:  coeff = 10'sd4; 
			9'd257:  coeff = 10'sd3; 
			9'd258:  coeff = 10'sd2; 
			9'd259:  coeff = 10'sd0; 
			9'd260:  coeff = -10'sd2; 
			9'd261:  coeff = -10'sd3; 
			9'd262:  coeff = -10'sd3; 
			9'd263:  coeff = -10'sd2; 
			9'd264:  coeff = -10'sd1; 
			9'd265:  coeff = 10'sd0; 
			9'd266:  coeff = 10'sd2; 
			9'd267:  coeff = 10'sd2; 
			9'd268:  coeff = 10'sd2; 
			9'd269:  coeff = 10'sd2; 
			9'd270:  coeff = 10'sd1; 
			9'd271:  coeff = 10'sd0; 
			9'd272:  coeff = -10'sd2; 
			9'd273:  coeff = -10'sd2; 
			9'd274:  coeff = -10'sd2; 
			9'd275:  coeff = -10'sd1; 
			9'd276:  coeff = 10'sd0; 
			9'd277:  coeff = 10'sd1; 
			9'd278:  coeff = 10'sd1; 
			9'd279:  coeff = 10'sd2; 
			9'd280:  coeff = 10'sd2; 
			9'd281:  coeff = 10'sd1; 
			9'd282:  coeff = 10'sd0; 
			9'd283:  coeff = -10'sd1; 
			9'd284:  coeff = -10'sd1; 
			9'd285:  coeff = -10'sd1; 
			9'd286:  coeff = -10'sd1; 
			9'd287:  coeff = -10'sd1; 
			9'd288:  coeff = 10'sd0; 
			9'd289:  coeff = 10'sd0; 
			9'd290:  coeff = 10'sd1; 
			9'd291:  coeff = 10'sd1; 
			9'd292:  coeff = 10'sd1; 
			9'd293:  coeff = 10'sd1; 
			9'd294:  coeff = 10'sd0; 
			9'd295:  coeff = 10'sd0; 
			9'd296:  coeff = -10'sd1; 
			9'd297:  coeff = -10'sd1; 
			9'd298:  coeff = -10'sd1; 
			9'd299:  coeff = 10'sd0; 
			9'd300:  coeff = 10'sd0; 
			9'd301:  coeff = 10'sd0; 
			9'd302:  coeff = 10'sd1; 
			9'd303:  coeff = 10'sd1; 
			9'd304:  coeff = 10'sd1; 
			9'd305:  coeff = 10'sd0; 
			9'd306:  coeff = 10'sd0; 
			9'd307:  coeff = 10'sd0; 
			9'd308:  coeff = -10'sd1; 
			9'd309:  coeff = -10'sd1; 
			9'd310:  coeff = 10'sd0; 
			9'd311:  coeff = 10'sd0; 
			9'd312:  coeff = 10'sd0; 
			9'd313:  coeff = 10'sd0; 
			9'd314:  coeff = 10'sd0; 
			9'd315:  coeff = 10'sd0; 
			9'd316:  coeff = 10'sd0; 
			9'd317:  coeff = 10'sd0; 
			9'd318:  coeff = 10'sd0; 
			9'd319:  coeff = 10'sd0; 
			9'd320:  coeff = 10'sd0; 
			9'd321:  coeff = 10'sd0; 
			9'd322:  coeff = 10'sd0; 
			9'd323:  coeff = 10'sd0; 
			9'd324:  coeff = 10'sd0; 
			9'd325:  coeff = 10'sd0; 
			9'd326:  coeff = 10'sd0; 
			9'd327:  coeff = 10'sd0; 
			9'd328:  coeff = 10'sd0; 
			9'd329:  coeff = 10'sd0; 
			9'd330:  coeff = 10'sd0; 
			9'd331:  coeff = 10'sd0; 
			9'd332:  coeff = 10'sd0; 
			9'd333:  coeff = 10'sd0; 
			9'd334:  coeff = 10'sd0; 
			9'd335:  coeff = 10'sd0; 
			9'd336:  coeff = 10'sd0; 
			9'd337:  coeff = 10'sd0; 
			9'd338:  coeff = 10'sd0; 
			9'd339:  coeff = 10'sd0; 
			9'd340:  coeff = 10'sd0; 
			9'd341:  coeff = 10'sd0; 
			9'd342:  coeff = 10'sd0; 
			9'd343:  coeff = 10'sd0; 
			9'd344:  coeff = 10'sd0; 
			9'd345:  coeff = 10'sd0; 
			9'd346:  coeff = 10'sd0; 
			9'd347:  coeff = 10'sd0; 
			9'd348:  coeff = 10'sd0; 
			9'd349:  coeff = 10'sd0; 
			9'd350:  coeff = 10'sd0; 
			9'd351:  coeff = 10'sd0; 
			9'd352:  coeff = 10'sd0; 
			9'd353:  coeff = 10'sd0; 
			9'd354:  coeff = 10'sd0; 
			9'd355:  coeff = 10'sd0; 
			9'd356:  coeff = 10'sd0; 
			9'd357:  coeff = 10'sd0; 
			9'd358:  coeff = 10'sd0; 
			9'd359:  coeff = 10'sd0; 
			9'd360:  coeff = 10'sd0; 
			9'd361:  coeff = 10'sd0; 
			9'd362:  coeff = 10'sd0; 
			9'd363:  coeff = 10'sd0; 
			9'd364:  coeff = 10'sd0; 
			9'd365:  coeff = 10'sd0; 
			9'd366:  coeff = 10'sd0; 
			9'd367:  coeff = 10'sd0; 
			9'd368:  coeff = 10'sd0; 
			9'd369:  coeff = 10'sd0; 
			9'd370:  coeff = 10'sd0; 
			9'd371:  coeff = 10'sd0; 
			9'd372:  coeff = 10'sd0; 
			9'd373:  coeff = 10'sd0; 
			9'd374:  coeff = 10'sd0; 
			9'd375:  coeff = 10'sd0; 
			9'd376:  coeff = 10'sd0; 
			9'd377:  coeff = 10'sd0; 
			9'd378:  coeff = 10'sd0; 
			9'd379:  coeff = 10'sd0; 
			9'd380:  coeff = 10'sd0; 
			9'd381:  coeff = 10'sd0; 
			9'd382:  coeff = 10'sd0; 
			9'd383:  coeff = 10'sd0; 
			9'd384:  coeff = 10'sd0; 
			9'd385:  coeff = 10'sd0; 
			9'd386:  coeff = 10'sd0; 
			9'd387:  coeff = 10'sd0; 
			9'd388:  coeff = 10'sd0; 
			9'd389:  coeff = 10'sd0; 
			9'd390:  coeff = 10'sd0; 
			9'd391:  coeff = 10'sd0; 
			9'd392:  coeff = 10'sd0; 
			9'd393:  coeff = 10'sd0; 
			9'd394:  coeff = 10'sd0; 
			9'd395:  coeff = 10'sd0; 
			9'd396:  coeff = 10'sd0; 
			9'd397:  coeff = 10'sd0; 
			9'd398:  coeff = 10'sd0; 
			9'd399:  coeff = 10'sd0; 
			9'd400:  coeff = 10'sd0; 

			default: coeff = 10'hXXX;
		endcase
endmodule

