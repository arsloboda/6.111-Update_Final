`default_nettype none

///////////////////////////////////////////////////////////////////////////////
//
// Switch Debounce Module
//
///////////////////////////////////////////////////////////////////////////////

module debounce (
  input wire reset, clock, noisy,
  output reg clean
);
  reg [18:0] count;
  reg new;

  always @(posedge clock)
    if (reset) begin
      count <= 0;
      new <= noisy;
      clean <= noisy;
    end
    else if (noisy != new) begin
      // noisy input changed, restart the .01 sec clock
      new <= noisy;
      count <= 0;
    end
    else if (count == 270000)
      // noisy input stable for .01 secs, pass it along!
      clean <= new;
    else
      // waiting for .01 sec to pass
      count <= count+1;

endmodule

///////////////////////////////////////////////////////////////////////////////
//
// bi-directional monaural 18bit interface to AC97
//
///////////////////////////////////////////////////////////////////////////////

module audio (
  input wire clock_27mhz,
  input wire reset,
  input wire [4:0] volume,
  output wire [17:0] left_audio_in_data,
  input wire [17:0] left_audio_out_data,
  output wire [17:0] right_audio_in_data,
  input wire [17:0] right_audio_out_data,
  output wire ready,
  output reg audio_reset_b,   // ac97 interface signals
  output wire ac97_sdata_out,
  input wire ac97_sdata_in,
  output wire ac97_synch,
  input wire ac97_bit_clock
);

  wire [7:0] command_address;
  wire [15:0] command_data;
  wire command_valid;
  wire [19:0] left_in_data, right_in_data;
  wire [19:0] left_out_data, right_out_data;

  // wait a little before enabling the AC97 codec
  reg [9:0] reset_count;
  always @(posedge clock_27mhz) begin
    if (reset) begin
      audio_reset_b = 1'b0;
      reset_count = 0;
    end else if (reset_count == 1023)
      audio_reset_b = 1'b1;
    else
      reset_count = reset_count+1;
  end

  wire ac97_ready;
  ac97 ac97(.ready(ac97_ready),
            .command_address(command_address),
            .command_data(command_data),
            .command_valid(command_valid),
            .left_data(left_out_data), .left_valid(1'b1),
            .right_data(right_out_data), .right_valid(1'b1),
            .left_in_data(left_in_data), .right_in_data(right_in_data),
            .ac97_sdata_out(ac97_sdata_out),
            .ac97_sdata_in(ac97_sdata_in),
            .ac97_synch(ac97_synch),
            .ac97_bit_clock(ac97_bit_clock));

  // ready: one cycle pulse synchronous with clock_27mhz
  reg [2:0] ready_sync;
  always @ (posedge clock_27mhz) ready_sync <= {ready_sync[1:0], ac97_ready};
  assign ready = ready_sync[1] & ~ready_sync[2];

  reg [17:0] out_data_l;
  reg [17:0] out_data_r;
  always @ (posedge clock_27mhz) begin
    if (ready) begin
		out_data_l <= left_audio_out_data;
		out_data_r <= right_audio_out_data;
	 end
  end
	 
  assign left_audio_in_data =  left_in_data[19:2];
  assign right_audio_in_data=  right_in_data[19:2];
  assign left_out_data ={out_data_l,2'b00};
  assign right_out_data={out_data_r,2'b00};

  // generate repeating sequence of read/writes to AC97 registers
  ac97commands cmds(.clock(clock_27mhz), .ready(ready),
                    .command_address(command_address),
                    .command_data(command_data),
                    .command_valid(command_valid),
                    .volume(volume),
                    .source(3'b100));     // mic
endmodule

// assemble/disassemble AC97 serial frames
module ac97 (
  output reg ready,
  input wire [7:0] command_address,
  input wire [15:0] command_data,
  input wire command_valid,
  input wire [19:0] left_data,
  input wire left_valid,
  input wire [19:0] right_data,
  input wire right_valid,
  output reg [19:0] left_in_data, right_in_data,
  output reg ac97_sdata_out,
  input wire ac97_sdata_in,
  output reg ac97_synch,
  input wire ac97_bit_clock
);
  reg [7:0] bit_count;

  reg [19:0] l_cmd_addr;
  reg [19:0] l_cmd_data;
  reg [19:0] l_left_data, l_right_data;
  reg l_cmd_v, l_left_v, l_right_v;

  initial begin
    ready <= 1'b0;
    // synthesis attribute init of ready is "0";
    ac97_sdata_out <= 1'b0;
    // synthesis attribute init of ac97_sdata_out is "0";
    ac97_synch <= 1'b0;
    // synthesis attribute init of ac97_synch is "0";

    bit_count <= 8'h00;
    // synthesis attribute init of bit_count is "0000";
    l_cmd_v <= 1'b0;
    // synthesis attribute init of l_cmd_v is "0";
    l_left_v <= 1'b0;
    // synthesis attribute init of l_left_v is "0";
    l_right_v <= 1'b0;
    // synthesis attribute init of l_right_v is "0";

    left_in_data <= 20'h00000;
    // synthesis attribute init of left_in_data is "00000";
    right_in_data <= 20'h00000;
    // synthesis attribute init of right_in_data is "00000";
  end

  always @(posedge ac97_bit_clock) begin
    // Generate the sync signal
    if (bit_count == 255)
      ac97_synch <= 1'b1;
    if (bit_count == 15)
      ac97_synch <= 1'b0;

    // Generate the ready signal
    if (bit_count == 128)
      ready <= 1'b1;
    if (bit_count == 2)
      ready <= 1'b0;

    // Latch user data at the end of each frame. This ensures that the
    // first frame after reset will be empty.
    if (bit_count == 255) begin
      l_cmd_addr <= {command_address, 12'h000};
      l_cmd_data <= {command_data, 4'h0};
      l_cmd_v <= command_valid;
      l_left_data <= left_data;
      l_left_v <= left_valid;
      l_right_data <= right_data;
      l_right_v <= right_valid;
    end

    if ((bit_count >= 0) && (bit_count <= 15))
      // Slot 0: Tags
      case (bit_count[3:0])
        4'h0: ac97_sdata_out <= 1'b1;      // Frame valid
        4'h1: ac97_sdata_out <= l_cmd_v;   // Command address valid
        4'h2: ac97_sdata_out <= l_cmd_v;   // Command data valid
        4'h3: ac97_sdata_out <= l_left_v;  // Left data valid
        4'h4: ac97_sdata_out <= l_right_v; // Right data valid
        default: ac97_sdata_out <= 1'b0;
      endcase
    else if ((bit_count >= 16) && (bit_count <= 35))
      // Slot 1: Command address (8-bits, left justified)
      ac97_sdata_out <= l_cmd_v ? l_cmd_addr[35-bit_count] : 1'b0;
    else if ((bit_count >= 36) && (bit_count <= 55))
      // Slot 2: Command data (16-bits, left justified)
      ac97_sdata_out <= l_cmd_v ? l_cmd_data[55-bit_count] : 1'b0;
    else if ((bit_count >= 56) && (bit_count <= 75)) begin
      // Slot 3: Left channel
      ac97_sdata_out <= l_left_v ? l_left_data[19] : 1'b0;
      l_left_data <= { l_left_data[18:0], l_left_data[19] };
    end
    else if ((bit_count >= 76) && (bit_count <= 95))
      // Slot 4: Right channel
      ac97_sdata_out <= l_right_v ? l_right_data[95-bit_count] : 1'b0;
    else
      ac97_sdata_out <= 1'b0;

    bit_count <= bit_count+1;
  end // always @ (posedge ac97_bit_clock)

  always @(negedge ac97_bit_clock) begin
    if ((bit_count >= 57) && (bit_count <= 76))
      // Slot 3: Left channel
      left_in_data <= { left_in_data[18:0], ac97_sdata_in };
    else if ((bit_count >= 77) && (bit_count <= 96))
      // Slot 4: Right channel
      right_in_data <= { right_in_data[18:0], ac97_sdata_in };
  end
endmodule

// issue initialization commands to AC97
module ac97commands (
  input wire clock,
  input wire ready,
  output wire [7:0] command_address,
  output wire [15:0] command_data,
  output reg command_valid,
  input wire [4:0] volume,
  input wire [2:0] source
);
  reg [23:0] command;

  reg [3:0] state;
  initial begin
    command <= 4'h0;
    // synthesis attribute init of command is "0";
    command_valid <= 1'b0;
    // synthesis attribute init of command_valid is "0";
    state <= 16'h0000;
    // synthesis attribute init of state is "0000";
  end

  assign command_address = command[23:16];
  assign command_data = command[15:0];

  wire [4:0] vol;
  assign vol = 31-volume;  // convert to attenuation

  always @(posedge clock) begin
    if (ready) state <= state+1;

    case (state)
      4'h0: // Read ID
        begin
          command <= 24'h80_0000;
          command_valid <= 1'b1;
        end
      4'h1: // Read ID
        command <= 24'h80_0000;
      4'h3: // headphone volume
        command <= { 8'h04, 3'b000, vol, 3'b000, vol };
      4'h5: // PCM volume
        command <= 24'h18_0808;
      4'h6: // Record source select
        command <= { 8'h1A, 5'b00000, source, 5'b00000, source};
      4'h7: // Record gain = max
        command <= 24'h1C_0F0F;
      4'h9: // set +20db mic gain
        command <= 24'h0E_8048;
      4'hA: // Set beep volume
        command <= 24'h0A_0000;
      4'hB: // PCM out bypass mix1
        command <= 24'h20_8000;
      default:
        command <= 24'h80_0000;
    endcase // case(state)
  end // always @ (posedge clock)
endmodule // ac97commands

/////////////////////////////////////////////////////////////////////////////////
////
//// 6.111 FPGA Labkit -- Template Toplevel Module
////
//// For Labkit Revision 004
//// Created: October 31, 2004, from revision 003 file
//// Author: Nathan Ickes, 6.111 staff
////
/////////////////////////////////////////////////////////////////////////////////

module Labkit_M   (beep, audio_reset_b, ac97_sdata_out, ac97_sdata_in, ac97_synch,
	       ac97_bit_clock,
	       
	       vga_out_red, vga_out_green, vga_out_blue, vga_out_sync_b,
	       vga_out_blank_b, vga_out_pixel_clock, vga_out_hsync,
	       vga_out_vsync,

	       tv_out_ycrcb, tv_out_reset_b, tv_out_clock, tv_out_i2c_clock,
	       tv_out_i2c_data, tv_out_pal_ntsc, tv_out_hsync_b,
	       tv_out_vsync_b, tv_out_blank_b, tv_out_subcar_reset,

	       tv_in_ycrcb, tv_in_data_valid, tv_in_line_clock1,
	       tv_in_line_clock2, tv_in_aef, tv_in_hff, tv_in_aff,
	       tv_in_i2c_clock, tv_in_i2c_data, tv_in_fifo_read,
	       tv_in_fifo_clock, tv_in_iso, tv_in_reset_b, tv_in_clock,

	       ram0_data, ram0_address, ram0_adv_ld, ram0_clk, ram0_cen_b,
	       ram0_ce_b, ram0_oe_b, ram0_we_b, ram0_bwe_b, 

	       ram1_data, ram1_address, ram1_adv_ld, ram1_clk, ram1_cen_b,
	       ram1_ce_b, ram1_oe_b, ram1_we_b, ram1_bwe_b,

	       clock_feedback_out, clock_feedback_in,

	       flash_data, flash_address, flash_ce_b, flash_oe_b, flash_we_b,
	       flash_reset_b, flash_sts, flash_byte_b,

	       rs232_txd, rs232_rxd, rs232_rts, rs232_cts,

	       mouse_clock, mouse_data, keyboard_clock, keyboard_data,

	       clock_27mhz, clock1, clock2,

	       disp_blank, disp_data_out, disp_clock, disp_rs, disp_ce_b,
	       disp_reset_b, disp_data_in,

	       button0, button1, button2, button3, button_enter, button_right,
	       button_left, button_down, button_up,

	       switch,

	       led,
	       
	       user1, user2, user3, user4,
	       
	       daughtercard,

	       systemace_data, systemace_address, systemace_ce_b,
	       systemace_we_b, systemace_oe_b, systemace_irq, systemace_mpbrdy,
	       
	       analyzer1_data, analyzer1_clock,
 	       analyzer2_data, analyzer2_clock,
 	       analyzer3_data, analyzer3_clock,
 	       analyzer4_data, analyzer4_clock);

   output beep, audio_reset_b, ac97_synch, ac97_sdata_out;
   input  ac97_bit_clock, ac97_sdata_in;
   
   output [7:0] vga_out_red, vga_out_green, vga_out_blue;
   output vga_out_sync_b, vga_out_blank_b, vga_out_pixel_clock,
	  vga_out_hsync, vga_out_vsync;

   output [9:0] tv_out_ycrcb;
   output tv_out_reset_b, tv_out_clock, tv_out_i2c_clock, tv_out_i2c_data,
	  tv_out_pal_ntsc, tv_out_hsync_b, tv_out_vsync_b, tv_out_blank_b,
	  tv_out_subcar_reset;
   
   input  [19:0] tv_in_ycrcb;
   input  tv_in_data_valid, tv_in_line_clock1, tv_in_line_clock2, tv_in_aef,
	  tv_in_hff, tv_in_aff;
   output tv_in_i2c_clock, tv_in_fifo_read, tv_in_fifo_clock, tv_in_iso,
	  tv_in_reset_b, tv_in_clock;
   inout  tv_in_i2c_data;
        
   inout  [35:0] ram0_data;
   output [18:0] ram0_address;
   output ram0_adv_ld, ram0_clk, ram0_cen_b, ram0_ce_b, ram0_oe_b, ram0_we_b;
   output [3:0] ram0_bwe_b;
   
   inout  [35:0] ram1_data;
   output [18:0] ram1_address;
   output ram1_adv_ld, ram1_clk, ram1_cen_b, ram1_ce_b, ram1_oe_b, ram1_we_b;
   output [3:0] ram1_bwe_b;

   input  clock_feedback_in;
   output clock_feedback_out;
   
   inout  [15:0] flash_data;
   output [23:0] flash_address;
   output flash_ce_b, flash_oe_b, flash_we_b, flash_reset_b, flash_byte_b;
   input  flash_sts;
   
   output rs232_txd, rs232_rts;
   input  rs232_rxd, rs232_cts;

   input  mouse_clock, mouse_data, keyboard_clock, keyboard_data;

   input  clock_27mhz, clock1, clock2;

   output disp_blank, disp_clock, disp_rs, disp_ce_b, disp_reset_b;  
   input  disp_data_in;
   output  disp_data_out;
   
   input  button0, button1, button2, button3, button_enter, button_right,
	  button_left, button_down, button_up;
   input  [7:0] switch;
   output [7:0] led;

   inout [31:0] user1, user2, user3, user4;
   
   inout [43:0] daughtercard;

   inout  [15:0] systemace_data;
   output [6:0]  systemace_address;
   output systemace_ce_b, systemace_we_b, systemace_oe_b;
   input  systemace_irq, systemace_mpbrdy;

   output [15:0] analyzer1_data, analyzer2_data, analyzer3_data, 
		 analyzer4_data;
   output analyzer1_clock, analyzer2_clock, analyzer3_clock, analyzer4_clock;

   ////////////////////////////////////////////////////////////////////////////
   //
   // I/O Assignments
   //
   ////////////////////////////////////////////////////////////////////////////
   

   // Audio Input and Output
   assign beep= 1'b0;
   //lab5 assign audio_reset_b = 1'b0;
   //lab5 assign ac97_synch = 1'b0;
   //lab5 assign ac97_sdata_out = 1'b0;
   // ac97_sdata_in is an input

   // VGA Output
   assign vga_out_red = 10'h0;
   assign vga_out_green = 10'h0;
   assign vga_out_blue = 10'h0;
   assign vga_out_sync_b = 1'b1;
   assign vga_out_blank_b = 1'b1;
   assign vga_out_pixel_clock = 1'b0;
   assign vga_out_hsync = 1'b0;
   assign vga_out_vsync = 1'b0;

   // Video Output
   assign tv_out_ycrcb = 10'h0;
   assign tv_out_reset_b = 1'b0;
   assign tv_out_clock = 1'b0;
   assign tv_out_i2c_clock = 1'b0;
   assign tv_out_i2c_data = 1'b0;
   assign tv_out_pal_ntsc = 1'b0;
   assign tv_out_hsync_b = 1'b1;
   assign tv_out_vsync_b = 1'b1;
   assign tv_out_blank_b = 1'b1;
   assign tv_out_subcar_reset = 1'b0;
   
   // Video Input
   assign tv_in_i2c_clock = 1'b0;
   assign tv_in_fifo_read = 1'b0;
   assign tv_in_fifo_clock = 1'b0;
   assign tv_in_iso = 1'b0;
   assign tv_in_reset_b = 1'b0;
   assign tv_in_clock = 1'b0;
   assign tv_in_i2c_data = 1'bZ;
   // tv_in_ycrcb, tv_in_data_valid, tv_in_line_clock1, tv_in_line_clock2, 
   // tv_in_aef, tv_in_hff, and tv_in_aff are inputs
   
   // SRAMs
   assign ram0_data = 36'hZ;
   assign ram0_address = 19'h0;
   assign ram0_adv_ld = 1'b0;
   assign ram0_clk = 1'b0;
   assign ram0_cen_b = 1'b1;
   assign ram0_ce_b = 1'b1;
   assign ram0_oe_b = 1'b1;
   assign ram0_we_b = 1'b1;
   assign ram0_bwe_b = 4'hF;
   assign ram1_data = 36'hZ; 
   assign ram1_address = 19'h0;
   assign ram1_adv_ld = 1'b0;
   assign ram1_clk = 1'b0;
   assign ram1_cen_b = 1'b1;
   assign ram1_ce_b = 1'b1;
   assign ram1_oe_b = 1'b1;
   assign ram1_we_b = 1'b1;
   assign ram1_bwe_b = 4'hF;
   assign clock_feedback_out = 1'b0;
   // clock_feedback_in is an input
   
//   // Flash ROM
//   assign flash_data = 16'hZ;
//   assign flash_address = 24'h0;
//   assign flash_ce_b = 1'b1;
//   assign flash_oe_b = 1'b1;
//   assign flash_we_b = 1'b1;
//   assign flash_reset_b = 1'b0;
//   assign flash_byte_b = 1'b1;
//   // flash_sts is an input

   // RS-232 Interface
   assign rs232_txd = 1'b1;
   assign rs232_rts = 1'b1;
   // rs232_rxd and rs232_cts are inputs

   // PS/2 Ports
   // mouse_clock, mouse_data, keyboard_clock, and keyboard_data are inputs

//   // LED Displays
//   assign disp_blank = 1'b1;
//   assign disp_clock = 1'b0;
//   assign disp_rs = 1'b0;
//   assign disp_ce_b = 1'b1;
//   assign disp_reset_b = 1'b0;
//   assign disp_data_out = 1'b0;
//   // disp_data_in is an input

   // Buttons, Switches, and Individual LEDs
   //lab5 assign led = 8'hFF;
   // button0, button1, button2, button3, button_enter, button_right,
   // button_left, button_down, button_up, and switches are inputs

   // User I/Os
   //assign user1 = 32'hZ;
   assign user2 = 32'hZ;
   assign user3 = 32'hZ;
//   assign user4 = 32'hZ;

   // Daughtercard Connectors
   assign daughtercard = 44'hZ;

   // SystemACE Microprocessor Port
   assign systemace_data = 16'hZ;
   assign systemace_address = 7'h0;
   assign systemace_ce_b = 1'b1;
   assign systemace_we_b = 1'b1;
   assign systemace_oe_b = 1'b1;
   // systemace_irq and systemace_mpbrdy are inputs

   // Logic Analyzer
   //lab5 assign analyzer1_data = 16'h0;
   //lab5 assign analyzer1_clock = 1'b1;
   assign analyzer2_data = 16'h0;
   assign analyzer2_clock = 1'b1;
   //lab5 assign analyzer3_data = 16'h0;
   //lab5 assign analyzer3_clock = 1'b1;
   assign analyzer4_data = 16'h0;
   assign analyzer4_clock = 1'b1;

   ////////////////////////////////////////////////////////////////////////////
   //
   // Reset Generation
   //
   // A shift register primitive is used to generate an active-high reset
   // signal that remains high for 16 clock cycles after configuration finishes
   // and the FPGA's internal clocks begin toggling.
   //
   ////////////////////////////////////////////////////////////////////////////
   wire reset;
   SRL16 #(.INIT(16'hFFFF)) reset_sr(.D(1'b0), .CLK(clock_27mhz), .Q(reset),
                                     .A0(1'b1), .A1(1'b1), .A2(1'b1), .A3(1'b1));

	////////////////////////////////////////////////////////////////////////////
	//
	// RELEVANT TOOLS FOR USING AUDIO INPUT AND OUTPUT
	//
	//
	//
	////////////////////////////////////////////////////////////////////////////
   wire [17:0] from_ac97_data_l, from_ac97_data_r;
   wire ready;
	
   // allow user to adjust volume
   wire vup,vdown,switch0,switch1,switch2,switch3,switch4;
	wire switch5,switch6,switch7,enter,reset2,b0,b1,b2,b3,bl,br;
   reg old_vup,old_vdown;
   debounce bup(.reset(reset),.clock(clock_27mhz),.noisy(~button_up),.clean(vup));
   debounce bdown(.reset(reset),.clock(clock_27mhz),.noisy(~button_down),.clean(vdown));
   debounce sw0(.reset(reset),.clock(clock_27mhz),.noisy(switch[0]),.clean(switch0));
   debounce sw1(.reset(reset),.clock(clock_27mhz),.noisy(switch[1]),.clean(switch1));
   debounce sw2(.reset(reset),.clock(clock_27mhz),.noisy(switch[2]),.clean(switch2));
	debounce sw3(.reset(reset),.clock(clock_27mhz),.noisy(switch[3]),.clean(switch3));
	debounce sw4(.reset(reset),.clock(clock_27mhz),.noisy(switch[4]),.clean(switch4));
	debounce sw5(.reset(reset),.clock(clock_27mhz),.noisy(switch[5]),.clean(switch5));
	debounce sw6(.reset(reset),.clock(clock_27mhz),.noisy(switch[6]),.clean(switch6));
	debounce sw7(.reset(reset),.clock(clock_27mhz),.noisy(switch[7]),.clean(switch7));
	debounce bent(.reset(reset),.clock(clock_27mhz),.noisy(~button_enter),.clean(enter));
   debounce but0(.reset(reset),.clock(clock_27mhz),.noisy(~button0),.clean(b0));
   debounce but1(.reset(reset),.clock(clock_27mhz),.noisy(~button1),.clean(b1));
   debounce but2(.reset(reset),.clock(clock_27mhz),.noisy(~button2),.clean(b2));
   debounce but3(.reset(reset),.clock(clock_27mhz),.noisy(~button3),.clean(b3));
   debounce butl(.reset(reset),.clock(clock_27mhz),.noisy(~button_left),.clean(bl));
   debounce butr(.reset(reset),.clock(clock_27mhz),.noisy(~button_right),.clean(br));

	reg [4:0] volume;
   always @ (posedge clock_27mhz) begin
     if (reset) volume <= 5'd24;
     else begin
	if (vup & ~old_vup & volume != 5'd31) volume <= volume+1;       
	if (vdown & ~old_vdown & volume != 5'd0) volume <= volume-1;       
     end
     old_vup <= vup;
     old_vdown <= vdown;
   end
	wire [17:0] for_ac97_l;
	wire [17:0] for_ac97_r;
	wire [9:0] f_controls;
	wire [9:0] t_controls;
	wire [9:0] m_controls;
	wire [11:0] status;
	wire [55:0] freq_data;
	
	// frequency weights output to hex display
	wire [4:0] test1;
	wire [4:0] test2;
	wire [4:0] test3;
	wire [4:0] test4;
	wire [4:0] test5;
	wire [4:0] test6;
	wire [4:0] test7;
	wire test_flash;
	wire test_flash2;
	wire do_record;
	wire do_play;
	wire writemode;
	
   //High Level FSM
	HighLevelFSM HLFSM(.clock(clock_27mhz),.reset(reset),
							.controls({bl,br,enter,b3,b2,b1,b0,switch7,
							switch6,switch5,switch4,switch3,switch2,switch1,switch0}),
							.f_controls(f_controls),.t_controls(t_controls),
							.m_controls(m_controls),
							.status(status));
	
	// AC97 driver
   audio a(clock_27mhz, reset, volume, from_ac97_data_l, for_ac97_l,from_ac97_data_r,for_ac97_r, ready,
	       audio_reset_b, ac97_sdata_out, ac97_sdata_in,
	       ac97_synch, ac97_bit_clock);
	
	//Assign output data
	ProcessMod process(.clock(clock_27mhz),.reset(reset),.ready(ready),
			 .l_audio_in(from_ac97_data_l),.r_audio_in(from_ac97_data_r),
			 .f_controls(f_controls),.t_controls(t_controls),
			 .l_audio_out(for_ac97_l),.r_audio_out(for_ac97_r),
			 .freq1(freq_data[7:0]),.freq2(freq_data[15:8]),
			 .freq3(freq_data[23:16]),.freq4(freq_data[31:24]),
			 .freq5(freq_data[39:32]),.freq6(freq_data[47:40]),
			 .freq7(freq_data[55:48]),.test1(test1),.test2(test2),
			 .test3(test3),.test4(test4),.test5(test5),.test6(test6),
			 .test7(test7));
			 
	wire [17:0] test_left;
	wire [17:0] test_right;	
	wire [15:0] frdata_check;
	music_flash_memory record_play(.clock(clock_27mhz),.reset(reset),.ready(ready),
//    		.do_record(do_record),.do_play(do_play),
				.left_audio_in(from_ac97_data_l),.right_audio_in(from_ac97_data_r),
				.flash_sts(flash_sts),.flash_data(flash_data),
//				.left_audio_out(for_ac97_l),.right_audio_out(for_ac97_r),
				.left_audio_out(test_left),.right_audio_out(test_right),
				.flash_address(flash_address),.flash_ce_b(flash_ce_b),
				.flash_oe_b(flash_oe_b),.flash_we_b(flash_we_b),
				.flash_reset_b(flash_reset_b),.flash_byte_b(flash_byte_b),
				.test(test_flash),.test2(test_flash2),
				.do_record(do_record),.do_play(do_play),.writemode(writemode),
				.frdata(frdata_check));
   
//	display_16hex disp(reset, clock_27mhz,
//			{240'b0,frdata_check}, // bits to output to hex display
//		
//			disp_blank, disp_clock, disp_rs, disp_ce_b,
//			disp_reset_b, disp_data_out);
	
	display_16hex disp(reset, clock_27mhz,
			{3'b0,test7,3'b0,test6,3'b0,test5,3'b0,test4,3'b0,test3,
			3'b0,test2,3'b0,test1}, // bits to output to hex display
		
			disp_blank, disp_clock, disp_rs, disp_ce_b,
			disp_reset_b, disp_data_out);
	
	
	wire [17:0] a_data;
   wire [29:0] LEDS;
	assign a_data=for_ac97_l;
	// show volume during playback.
   // led is active low
   assign led = ~{status[11:10],switch0, volume};
//   assign led = ~{writemode,do_record,do_play, volume};
   VDM lights(.clock(clock_27mhz),.reset(reset),.ready(ready),
              .a_data(a_data[17:0]),.f_data(48'b0),.controls(1'b0),
              .lights(LEDS));

   assign user4[4:0]=~{LEDS[4:0]};
   assign user4[12:8]=~{LEDS[9:5]};
   assign user4[20:16]=~{LEDS[14:10]};
   assign user3[4:0]=~{LEDS[19:15]};
   assign user3[12:8]=~{LEDS[24:20]};
   assign user3[20:16]=~{LEDS[29:25]};
   // output useful things to the logic analyzer connectors
   assign analyzer1_clock = ac97_bit_clock;
   assign analyzer1_data[0] = audio_reset_b;
   assign analyzer1_data[1] = ac97_sdata_out;
   assign analyzer1_data[2] = ac97_sdata_in;
   assign analyzer1_data[3] = ac97_synch;
   assign analyzer1_data[15:4] = 0;

   assign analyzer3_clock = ready;
   assign analyzer3_data = {from_ac97_data_l, for_ac97_l};
endmodule

///////////////////////////////////////////////////////////////////////////////
/// Hex Display Module
///////////////////////////////////////////////////////////////////////////////

module display_16hex (reset, clock_27mhz, data, 
		disp_blank, disp_clock, disp_rs, disp_ce_b,
		disp_reset_b, disp_data_out);

   input reset, clock_27mhz;    // clock and reset (active high reset)
   input [63:0] data;		// 16 hex nibbles to display
   
   output disp_blank, disp_clock, disp_data_out, disp_rs, disp_ce_b, 
	  disp_reset_b;
   
   reg disp_data_out, disp_rs, disp_ce_b, disp_reset_b;
   
   ////////////////////////////////////////////////////////////////////////////
   //
   // Display Clock
   //
   // Generate a 500kHz clock for driving the displays.
   //
   ////////////////////////////////////////////////////////////////////////////
   
   reg [4:0] count;
   reg [7:0] reset_count;
   reg clock;
   wire dreset;

   always @(posedge clock_27mhz)
     begin
	if (reset)
	  begin
	     count = 0;
	     clock = 0;
	  end
	else if (count == 26)
	  begin
	     clock = ~clock;
	     count = 5'h00;
	  end
	else
	  count = count+1;
     end
   
   always @(posedge clock_27mhz)
     if (reset)
       reset_count <= 100;
     else
       reset_count <= (reset_count==0) ? 0 : reset_count-1;

   assign dreset = (reset_count != 0);

   assign disp_clock = ~clock;

   ////////////////////////////////////////////////////////////////////////////
   //
   // Display State Machine
   //
   ////////////////////////////////////////////////////////////////////////////
      
   reg [7:0] state;		// FSM state
   reg [9:0] dot_index;		// index to current dot being clocked out
   reg [31:0] control;		// control register
   reg [3:0] char_index;	// index of current character
   reg [39:0] dots;		// dots for a single digit 
   reg [3:0] nibble;		// hex nibble of current character
   
   assign disp_blank = 1'b0; // low <= not blanked
   
   always @(posedge clock)
     if (dreset)
       begin
	  state <= 0;
	  dot_index <= 0;
	  control <= 32'h7F7F7F7F;
       end
     else
       casex (state)
	 8'h00:
	   begin
	      // Reset displays
	      disp_data_out <= 1'b0; 
	      disp_rs <= 1'b0; // dot register
	      disp_ce_b <= 1'b1;
	      disp_reset_b <= 1'b0;	     
	      dot_index <= 0;
	      state <= state+1;
	   end
	 
	 8'h01:
	   begin
	      // End reset
	      disp_reset_b <= 1'b1;
	      state <= state+1;
	   end
	 
	 8'h02:
	   begin
	      // Initialize dot register (set all dots to zero)
	      disp_ce_b <= 1'b0;
	      disp_data_out <= 1'b0; // dot_index[0];
	      if (dot_index == 639)
		state <= state+1;
	      else
		dot_index <= dot_index+1;
	   end
	 
	 8'h03:
	   begin
	      // Latch dot data
	      disp_ce_b <= 1'b1;
	      dot_index <= 31;		// re-purpose to init ctrl reg
	      disp_rs <= 1'b1; // Select the control register
	      state <= state+1;
	   end
	 
	 8'h04:
	   begin
	      // Setup the control register
	      disp_ce_b <= 1'b0;
	      disp_data_out <= control[31];
	      control <= {control[30:0], 1'b0};	// shift left
	      if (dot_index == 0)
		state <= state+1;
	      else
		dot_index <= dot_index-1;
	   end
	  
	 8'h05:
	   begin
	      // Latch the control register data / dot data
	      disp_ce_b <= 1'b1;
	      dot_index <= 39;		// init for single char
	      char_index <= 15;		// start with MS char
	      state <= state+1;
	      disp_rs <= 1'b0;	 	// Select the dot register
	   end
	 
	 8'h06:
	   begin
	      // Load the user's dot data into the dot reg, char by char
	      disp_ce_b <= 1'b0;
	      disp_data_out <= dots[dot_index]; // dot data from msb
	      if (dot_index == 0)
	        if (char_index == 0)
	          state <= 5;			// all done, latch data
		else
		begin
		  char_index <= char_index - 1;	// goto next char
		  dot_index <= 39;
		end
	      else
		dot_index <= dot_index-1;	// else loop thru all dots 
	   end

       endcase

   always @ (data or char_index)
     case (char_index)
       4'h0: 	 	nibble <= data[3:0];
       4'h1: 	 	nibble <= data[7:4];
       4'h2: 	 	nibble <= data[11:8];
       4'h3: 	 	nibble <= data[15:12];
       4'h4: 	 	nibble <= data[19:16];
       4'h5: 	 	nibble <= data[23:20];
       4'h6: 	 	nibble <= data[27:24];
       4'h7: 	 	nibble <= data[31:28];
       4'h8: 	 	nibble <= data[35:32];
       4'h9: 	 	nibble <= data[39:36];
       4'hA: 	 	nibble <= data[43:40];
       4'hB: 	 	nibble <= data[47:44];
       4'hC: 	 	nibble <= data[51:48];
       4'hD: 	 	nibble <= data[55:52];
       4'hE: 	 	nibble <= data[59:56];
       4'hF: 	 	nibble <= data[63:60];
     endcase
      
   always @(nibble)
     case (nibble)
       4'h0: dots <= 40'b00111110_01010001_01001001_01000101_00111110;
       4'h1: dots <= 40'b00000000_01000010_01111111_01000000_00000000;
       4'h2: dots <= 40'b01100010_01010001_01001001_01001001_01000110;
       4'h3: dots <= 40'b00100010_01000001_01001001_01001001_00110110;
       4'h4: dots <= 40'b00011000_00010100_00010010_01111111_00010000;
       4'h5: dots <= 40'b00100111_01000101_01000101_01000101_00111001;
       4'h6: dots <= 40'b00111100_01001010_01001001_01001001_00110000;
       4'h7: dots <= 40'b00000001_01110001_00001001_00000101_00000011;
       4'h8: dots <= 40'b00110110_01001001_01001001_01001001_00110110;
       4'h9: dots <= 40'b00000110_01001001_01001001_00101001_00011110;
       4'hA: dots <= 40'b01111110_00001001_00001001_00001001_01111110;
       4'hB: dots <= 40'b01111111_01001001_01001001_01001001_00110110;
       4'hC: dots <= 40'b00111110_01000001_01000001_01000001_00100010;
       4'hD: dots <= 40'b01111111_01000001_01000001_01000001_00111110;
       4'hE: dots <= 40'b01111111_01001001_01001001_01001001_01000001;
       4'hF: dots <= 40'b01111111_00001001_00001001_00001001_00000001;
     endcase
   
endmodule













//`default_nettype none
//
/////////////////////////////////////////////////////////////////////////////////
////
//// Switch Debounce Module
////
/////////////////////////////////////////////////////////////////////////////////
//
//module debounce (
//  input wire reset, clock, noisy,
//  output reg clean
//);
//  reg [18:0] count;
//  reg new;
//
//  always @(posedge clock)
//    if (reset) begin
//      count <= 0;
//      new <= noisy;
//      clean <= noisy;
//    end
//    else if (noisy != new) begin
//      // noisy input changed, restart the .01 sec clock
//      new <= noisy;
//      count <= 0;
//    end
//    else if (count == 270000)
//      // noisy input stable for .01 secs, pass it along!
//      clean <= new;
//    else
//      // waiting for .01 sec to pass
//      count <= count+1;
//
//endmodule
//
/////////////////////////////////////////////////////////////////////////////////
////
//// bi-directional monaural 18bit interface to AC97
////
/////////////////////////////////////////////////////////////////////////////////
//
//module audio (
//  input wire clock_27mhz,
//  input wire reset,
//  input wire [4:0] volume,
//  output wire [17:0] left_audio_in_data,
//  input wire [17:0] left_audio_out_data,
//  output wire [17:0] right_audio_in_data,
//  input wire [17:0] right_audio_out_data,
//  output wire ready,
//  output reg audio_reset_b,   // ac97 interface signals
//  output wire ac97_sdata_out,
//  input wire ac97_sdata_in,
//  output wire ac97_synch,
//  input wire ac97_bit_clock
//);
//
//  wire [7:0] command_address;
//  wire [15:0] command_data;
//  wire command_valid;
//  wire [19:0] left_in_data, right_in_data;
//  wire [19:0] left_out_data, right_out_data;
//
//  // wait a little before enabling the AC97 codec
//  reg [9:0] reset_count;
//  always @(posedge clock_27mhz) begin
//    if (reset) begin
//      audio_reset_b = 1'b0;
//      reset_count = 0;
//    end else if (reset_count == 1023)
//      audio_reset_b = 1'b1;
//    else
//      reset_count = reset_count+1;
//  end
//
//  wire ac97_ready;
//  ac97 ac97(.ready(ac97_ready),
//            .command_address(command_address),
//            .command_data(command_data),
//            .command_valid(command_valid),
//            .left_data(left_out_data), .left_valid(1'b1),
//            .right_data(right_out_data), .right_valid(1'b1),
//            .left_in_data(left_in_data), .right_in_data(right_in_data),
//            .ac97_sdata_out(ac97_sdata_out),
//            .ac97_sdata_in(ac97_sdata_in),
//            .ac97_synch(ac97_synch),
//            .ac97_bit_clock(ac97_bit_clock));
//
//  // ready: one cycle pulse synchronous with clock_27mhz
//  reg [2:0] ready_sync;
//  always @ (posedge clock_27mhz) ready_sync <= {ready_sync[1:0], ac97_ready};
//  assign ready = ready_sync[1] & ~ready_sync[2];
//
//  reg [17:0] out_data_l;
//  reg [17:0] out_data_r;
//  always @ (posedge clock_27mhz) begin
//    if (ready) begin
//		out_data_l <= left_audio_out_data;
//		out_data_r <= right_audio_out_data;
//	 end
//  end
//	 
//  assign left_audio_in_data =  left_in_data[19:2];
//  assign right_audio_in_data=  right_in_data[19:2];
//  assign left_out_data ={out_data_l,2'b00};
//  assign right_out_data={out_data_r,2'b00};
//
//  // generate repeating sequence of read/writes to AC97 registers
//  ac97commands cmds(.clock(clock_27mhz), .ready(ready),
//                    .command_address(command_address),
//                    .command_data(command_data),
//                    .command_valid(command_valid),
//                    .volume(volume),
//                    .source(3'b100));     // mic
//endmodule
//
//// assemble/disassemble AC97 serial frames
//module ac97 (
//  output reg ready,
//  input wire [7:0] command_address,
//  input wire [15:0] command_data,
//  input wire command_valid,
//  input wire [19:0] left_data,
//  input wire left_valid,
//  input wire [19:0] right_data,
//  input wire right_valid,
//  output reg [19:0] left_in_data, right_in_data,
//  output reg ac97_sdata_out,
//  input wire ac97_sdata_in,
//  output reg ac97_synch,
//  input wire ac97_bit_clock
//);
//  reg [7:0] bit_count;
//
//  reg [19:0] l_cmd_addr;
//  reg [19:0] l_cmd_data;
//  reg [19:0] l_left_data, l_right_data;
//  reg l_cmd_v, l_left_v, l_right_v;
//
//  initial begin
//    ready <= 1'b0;
//    // synthesis attribute init of ready is "0";
//    ac97_sdata_out <= 1'b0;
//    // synthesis attribute init of ac97_sdata_out is "0";
//    ac97_synch <= 1'b0;
//    // synthesis attribute init of ac97_synch is "0";
//
//    bit_count <= 8'h00;
//    // synthesis attribute init of bit_count is "0000";
//    l_cmd_v <= 1'b0;
//    // synthesis attribute init of l_cmd_v is "0";
//    l_left_v <= 1'b0;
//    // synthesis attribute init of l_left_v is "0";
//    l_right_v <= 1'b0;
//    // synthesis attribute init of l_right_v is "0";
//
//    left_in_data <= 20'h00000;
//    // synthesis attribute init of left_in_data is "00000";
//    right_in_data <= 20'h00000;
//    // synthesis attribute init of right_in_data is "00000";
//  end
//
//  always @(posedge ac97_bit_clock) begin
//    // Generate the sync signal
//    if (bit_count == 255)
//      ac97_synch <= 1'b1;
//    if (bit_count == 15)
//      ac97_synch <= 1'b0;
//
//    // Generate the ready signal
//    if (bit_count == 128)
//      ready <= 1'b1;
//    if (bit_count == 2)
//      ready <= 1'b0;
//
//    // Latch user data at the end of each frame. This ensures that the
//    // first frame after reset will be empty.
//    if (bit_count == 255) begin
//      l_cmd_addr <= {command_address, 12'h000};
//      l_cmd_data <= {command_data, 4'h0};
//      l_cmd_v <= command_valid;
//      l_left_data <= left_data;
//      l_left_v <= left_valid;
//      l_right_data <= right_data;
//      l_right_v <= right_valid;
//    end
//
//    if ((bit_count >= 0) && (bit_count <= 15))
//      // Slot 0: Tags
//      case (bit_count[3:0])
//        4'h0: ac97_sdata_out <= 1'b1;      // Frame valid
//        4'h1: ac97_sdata_out <= l_cmd_v;   // Command address valid
//        4'h2: ac97_sdata_out <= l_cmd_v;   // Command data valid
//        4'h3: ac97_sdata_out <= l_left_v;  // Left data valid
//        4'h4: ac97_sdata_out <= l_right_v; // Right data valid
//        default: ac97_sdata_out <= 1'b0;
//      endcase
//    else if ((bit_count >= 16) && (bit_count <= 35))
//      // Slot 1: Command address (8-bits, left justified)
//      ac97_sdata_out <= l_cmd_v ? l_cmd_addr[35-bit_count] : 1'b0;
//    else if ((bit_count >= 36) && (bit_count <= 55))
//      // Slot 2: Command data (16-bits, left justified)
//      ac97_sdata_out <= l_cmd_v ? l_cmd_data[55-bit_count] : 1'b0;
//    else if ((bit_count >= 56) && (bit_count <= 75)) begin
//      // Slot 3: Left channel
//      ac97_sdata_out <= l_left_v ? l_left_data[19] : 1'b0;
//      l_left_data <= { l_left_data[18:0], l_left_data[19] };
//    end
//    else if ((bit_count >= 76) && (bit_count <= 95))
//      // Slot 4: Right channel
//      ac97_sdata_out <= l_right_v ? l_right_data[95-bit_count] : 1'b0;
//    else
//      ac97_sdata_out <= 1'b0;
//
//    bit_count <= bit_count+1;
//  end // always @ (posedge ac97_bit_clock)
//
//  always @(negedge ac97_bit_clock) begin
//    if ((bit_count >= 57) && (bit_count <= 76))
//      // Slot 3: Left channel
//      left_in_data <= { left_in_data[18:0], ac97_sdata_in };
//    else if ((bit_count >= 77) && (bit_count <= 96))
//      // Slot 4: Right channel
//      right_in_data <= { right_in_data[18:0], ac97_sdata_in };
//  end
//endmodule
//
//// issue initialization commands to AC97
//module ac97commands (
//  input wire clock,
//  input wire ready,
//  output wire [7:0] command_address,
//  output wire [15:0] command_data,
//  output reg command_valid,
//  input wire [4:0] volume,
//  input wire [2:0] source
//);
//  reg [23:0] command;
//
//  reg [3:0] state;
//  initial begin
//    command <= 4'h0;
//    // synthesis attribute init of command is "0";
//    command_valid <= 1'b0;
//    // synthesis attribute init of command_valid is "0";
//    state <= 16'h0000;
//    // synthesis attribute init of state is "0000";
//  end
//
//  assign command_address = command[23:16];
//  assign command_data = command[15:0];
//
//  wire [4:0] vol;
//  assign vol = 31-volume;  // convert to attenuation
//
//  always @(posedge clock) begin
//    if (ready) state <= state+1;
//
//    case (state)
//      4'h0: // Read ID
//        begin
//          command <= 24'h80_0000;
//          command_valid <= 1'b1;
//        end
//      4'h1: // Read ID
//        command <= 24'h80_0000;
//      4'h3: // headphone volume
//        command <= { 8'h04, 3'b000, vol, 3'b000, vol };
//      4'h5: // PCM volume
//        command <= 24'h18_0808;
//      4'h6: // Record source select
//        command <= { 8'h1A, 5'b00000, source, 5'b00000, source};
//      4'h7: // Record gain = max
//        command <= 24'h1C_0F0F;
//      4'h9: // set +20db mic gain
//        command <= 24'h0E_8048;
//      4'hA: // Set beep volume
//        command <= 24'h0A_0000;
//      4'hB: // PCM out bypass mix1
//        command <= 24'h20_8000;
//      default:
//        command <= 24'h80_0000;
//    endcase // case(state)
//  end // always @ (posedge clock)
//endmodule // ac97commands
//
///////////////////////////////////////////////////////////////////////////////////
//////
////// 6.111 FPGA Labkit -- Template Toplevel Module
//////
////// For Labkit Revision 004
////// Created: October 31, 2004, from revision 003 file
////// Author: Nathan Ickes, 6.111 staff
//////
///////////////////////////////////////////////////////////////////////////////////
//
//module Labkit_M   (beep, audio_reset_b, ac97_sdata_out, ac97_sdata_in, ac97_synch,
//	       ac97_bit_clock,
//	       
//	       vga_out_red, vga_out_green, vga_out_blue, vga_out_sync_b,
//	       vga_out_blank_b, vga_out_pixel_clock, vga_out_hsync,
//	       vga_out_vsync,
//
//	       tv_out_ycrcb, tv_out_reset_b, tv_out_clock, tv_out_i2c_clock,
//	       tv_out_i2c_data, tv_out_pal_ntsc, tv_out_hsync_b,
//	       tv_out_vsync_b, tv_out_blank_b, tv_out_subcar_reset,
//
//	       tv_in_ycrcb, tv_in_data_valid, tv_in_line_clock1,
//	       tv_in_line_clock2, tv_in_aef, tv_in_hff, tv_in_aff,
//	       tv_in_i2c_clock, tv_in_i2c_data, tv_in_fifo_read,
//	       tv_in_fifo_clock, tv_in_iso, tv_in_reset_b, tv_in_clock,
//
//	       ram0_data, ram0_address, ram0_adv_ld, ram0_clk, ram0_cen_b,
//	       ram0_ce_b, ram0_oe_b, ram0_we_b, ram0_bwe_b, 
//
//	       ram1_data, ram1_address, ram1_adv_ld, ram1_clk, ram1_cen_b,
//	       ram1_ce_b, ram1_oe_b, ram1_we_b, ram1_bwe_b,
//
//	       clock_feedback_out, clock_feedback_in,
//
//	       flash_data, flash_address, flash_ce_b, flash_oe_b, flash_we_b,
//	       flash_reset_b, flash_sts, flash_byte_b,
//
//	       rs232_txd, rs232_rxd, rs232_rts, rs232_cts,
//
//	       mouse_clock, mouse_data, keyboard_clock, keyboard_data,
//
//	       clock_27mhz, clock1, clock2,
//
//	       disp_blank, disp_data_out, disp_clock, disp_rs, disp_ce_b,
//	       disp_reset_b, disp_data_in,
//
//	       button0, button1, button2, button3, button_enter, button_right,
//	       button_left, button_down, button_up,
//
//	       switch,
//
//	       led,
//	       
//	       user1, user2, user3, user4,
//	       
//	       daughtercard,
//
//	       systemace_data, systemace_address, systemace_ce_b,
//	       systemace_we_b, systemace_oe_b, systemace_irq, systemace_mpbrdy,
//	       
//	       analyzer1_data, analyzer1_clock,
// 	       analyzer2_data, analyzer2_clock,
// 	       analyzer3_data, analyzer3_clock,
// 	       analyzer4_data, analyzer4_clock);
//
//   output beep, audio_reset_b, ac97_synch, ac97_sdata_out;
//   input  ac97_bit_clock, ac97_sdata_in;
//   
//   output [7:0] vga_out_red, vga_out_green, vga_out_blue;
//   output vga_out_sync_b, vga_out_blank_b, vga_out_pixel_clock,
//	  vga_out_hsync, vga_out_vsync;
//
//   output [9:0] tv_out_ycrcb;
//   output tv_out_reset_b, tv_out_clock, tv_out_i2c_clock, tv_out_i2c_data,
//	  tv_out_pal_ntsc, tv_out_hsync_b, tv_out_vsync_b, tv_out_blank_b,
//	  tv_out_subcar_reset;
//   
//   input  [19:0] tv_in_ycrcb;
//   input  tv_in_data_valid, tv_in_line_clock1, tv_in_line_clock2, tv_in_aef,
//	  tv_in_hff, tv_in_aff;
//   output tv_in_i2c_clock, tv_in_fifo_read, tv_in_fifo_clock, tv_in_iso,
//	  tv_in_reset_b, tv_in_clock;
//   inout  tv_in_i2c_data;
//        
//   inout  [35:0] ram0_data;
//   output [18:0] ram0_address;
//   output ram0_adv_ld, ram0_clk, ram0_cen_b, ram0_ce_b, ram0_oe_b, ram0_we_b;
//   output [3:0] ram0_bwe_b;
//   
//   inout  [35:0] ram1_data;
//   output [18:0] ram1_address;
//   output ram1_adv_ld, ram1_clk, ram1_cen_b, ram1_ce_b, ram1_oe_b, ram1_we_b;
//   output [3:0] ram1_bwe_b;
//
//   input  clock_feedback_in;
//   output clock_feedback_out;
//   
//   inout  [15:0] flash_data;
//   output [23:0] flash_address;
//   output flash_ce_b, flash_oe_b, flash_we_b, flash_reset_b, flash_byte_b;
//   input  flash_sts;
//   
//   output rs232_txd, rs232_rts;
//   input  rs232_rxd, rs232_cts;
//
//   input  mouse_clock, mouse_data, keyboard_clock, keyboard_data;
//
//   input  clock_27mhz, clock1, clock2;
//
//   output disp_blank, disp_clock, disp_rs, disp_ce_b, disp_reset_b;  
//   input  disp_data_in;
//   output  disp_data_out;
//   
//   input  button0, button1, button2, button3, button_enter, button_right,
//	  button_left, button_down, button_up;
//   input  [7:0] switch;
//   output [7:0] led;
//
//   inout [31:0] user1, user2, user3, user4;
//   
//   inout [43:0] daughtercard;
//
//   inout  [15:0] systemace_data;
//   output [6:0]  systemace_address;
//   output systemace_ce_b, systemace_we_b, systemace_oe_b;
//   input  systemace_irq, systemace_mpbrdy;
//
//   output [15:0] analyzer1_data, analyzer2_data, analyzer3_data, 
//		 analyzer4_data;
//   output analyzer1_clock, analyzer2_clock, analyzer3_clock, analyzer4_clock;
//
//   ////////////////////////////////////////////////////////////////////////////
//   //
//   // I/O Assignments
//   //
//   ////////////////////////////////////////////////////////////////////////////
//   
//
//   // Audio Input and Output
//   assign beep= 1'b0;
//   //lab5 assign audio_reset_b = 1'b0;
//   //lab5 assign ac97_synch = 1'b0;
//   //lab5 assign ac97_sdata_out = 1'b0;
//   // ac97_sdata_in is an input
//
//   // VGA Output
//   assign vga_out_red = 10'h0;
//   assign vga_out_green = 10'h0;
//   assign vga_out_blue = 10'h0;
//   assign vga_out_sync_b = 1'b1;
//   assign vga_out_blank_b = 1'b1;
//   assign vga_out_pixel_clock = 1'b0;
//   assign vga_out_hsync = 1'b0;
//   assign vga_out_vsync = 1'b0;
//
//   // Video Output
//   assign tv_out_ycrcb = 10'h0;
//   assign tv_out_reset_b = 1'b0;
//   assign tv_out_clock = 1'b0;
//   assign tv_out_i2c_clock = 1'b0;
//   assign tv_out_i2c_data = 1'b0;
//   assign tv_out_pal_ntsc = 1'b0;
//   assign tv_out_hsync_b = 1'b1;
//   assign tv_out_vsync_b = 1'b1;
//   assign tv_out_blank_b = 1'b1;
//   assign tv_out_subcar_reset = 1'b0;
//   
//   // Video Input
//   assign tv_in_i2c_clock = 1'b0;
//   assign tv_in_fifo_read = 1'b0;
//   assign tv_in_fifo_clock = 1'b0;
//   assign tv_in_iso = 1'b0;
//   assign tv_in_reset_b = 1'b0;
//   assign tv_in_clock = 1'b0;
//   assign tv_in_i2c_data = 1'bZ;
//   // tv_in_ycrcb, tv_in_data_valid, tv_in_line_clock1, tv_in_line_clock2, 
//   // tv_in_aef, tv_in_hff, and tv_in_aff are inputs
//   
//   // SRAMs
//   assign ram0_data = 36'hZ;
//   assign ram0_address = 19'h0;
//   assign ram0_adv_ld = 1'b0;
//   assign ram0_clk = 1'b0;
//   assign ram0_cen_b = 1'b1;
//   assign ram0_ce_b = 1'b1;
//   assign ram0_oe_b = 1'b1;
//   assign ram0_we_b = 1'b1;
//   assign ram0_bwe_b = 4'hF;
//   assign ram1_data = 36'hZ; 
//   assign ram1_address = 19'h0;
//   assign ram1_adv_ld = 1'b0;
//   assign ram1_clk = 1'b0;
//   assign ram1_cen_b = 1'b1;
//   assign ram1_ce_b = 1'b1;
//   assign ram1_oe_b = 1'b1;
//   assign ram1_we_b = 1'b1;
//   assign ram1_bwe_b = 4'hF;
//   assign clock_feedback_out = 1'b0;
//   // clock_feedback_in is an input
//   
//   // Flash ROM
//   assign flash_data = 16'hZ;
//   assign flash_address = 24'h0;
//   assign flash_ce_b = 1'b1;
//   assign flash_oe_b = 1'b1;
//   assign flash_we_b = 1'b1;
//   assign flash_reset_b = 1'b0;
//   assign flash_byte_b = 1'b1;
//   // flash_sts is an input
//
//   // RS-232 Interface
//   assign rs232_txd = 1'b1;
//   assign rs232_rts = 1'b1;
//   // rs232_rxd and rs232_cts are inputs
//
//   // PS/2 Ports
//   // mouse_clock, mouse_data, keyboard_clock, and keyboard_data are inputs
//
////   // LED Displays
////   assign disp_blank = 1'b1;
////   assign disp_clock = 1'b0;
////   assign disp_rs = 1'b0;
////   assign disp_ce_b = 1'b1;
////   assign disp_reset_b = 1'b0;
////   assign disp_data_out = 1'b0;
////   // disp_data_in is an input
//
//   // Buttons, Switches, and Individual LEDs
//   //lab5 assign led = 8'hFF;
//   // button0, button1, button2, button3, button_enter, button_right,
//   // button_left, button_down, button_up, and switches are inputs
//
//   // User I/Os
//   //assign user1 = 32'hZ;
//   assign user2 = 32'hZ;
//   assign user3 = 32'hZ;
////   assign user4 = 32'hZ;
//
//   // Daughtercard Connectors
//   assign daughtercard = 44'hZ;
//
//   // SystemACE Microprocessor Port
//   assign systemace_data = 16'hZ;
//   assign systemace_address = 7'h0;
//   assign systemace_ce_b = 1'b1;
//   assign systemace_we_b = 1'b1;
//   assign systemace_oe_b = 1'b1;
//   // systemace_irq and systemace_mpbrdy are inputs
//
//   // Logic Analyzer
//   //lab5 assign analyzer1_data = 16'h0;
//   //lab5 assign analyzer1_clock = 1'b1;
//   assign analyzer2_data = 16'h0;
//   assign analyzer2_clock = 1'b1;
//   //lab5 assign analyzer3_data = 16'h0;
//   //lab5 assign analyzer3_clock = 1'b1;
//   assign analyzer4_data = 16'h0;
//   assign analyzer4_clock = 1'b1;
//
//   ////////////////////////////////////////////////////////////////////////////
//   //
//   // Reset Generation
//   //
//   // A shift register primitive is used to generate an active-high reset
//   // signal that remains high for 16 clock cycles after configuration finishes
//   // and the FPGA's internal clocks begin toggling.
//   //
//   ////////////////////////////////////////////////////////////////////////////
//   wire reset;
//   SRL16 #(.INIT(16'hFFFF)) reset_sr(.D(1'b0), .CLK(clock_27mhz), .Q(reset),
//                                     .A0(1'b1), .A1(1'b1), .A2(1'b1), .A3(1'b1));
//
//	////////////////////////////////////////////////////////////////////////////
//	//
//	// RELEVANT TOOLS FOR USING AUDIO INPUT AND OUTPUT
//	//
//	//
//	//
//	////////////////////////////////////////////////////////////////////////////
//   wire [17:0] from_ac97_data_l, from_ac97_data_r;
//   wire ready;
//	
//   // allow user to adjust volume
//   wire vup,vdown,switch0,switch1,switch2,switch3,switch4;
//	wire switch5,switch6,switch7,enter,reset2,b0,b1,b2,b3,bl,br;
//   reg old_vup,old_vdown;
//   debounce bup(.reset(reset),.clock(clock_27mhz),.noisy(~button_up),.clean(vup));
//   debounce bdown(.reset(reset),.clock(clock_27mhz),.noisy(~button_down),.clean(vdown));
//   debounce sw0(.reset(reset),.clock(clock_27mhz),.noisy(switch[0]),.clean(switch0));
//   debounce sw1(.reset(reset),.clock(clock_27mhz),.noisy(switch[1]),.clean(switch1));
//   debounce sw2(.reset(reset),.clock(clock_27mhz),.noisy(switch[2]),.clean(switch2));
//	debounce sw3(.reset(reset),.clock(clock_27mhz),.noisy(switch[3]),.clean(switch3));
//	debounce sw4(.reset(reset),.clock(clock_27mhz),.noisy(switch[4]),.clean(switch4));
//	debounce sw5(.reset(reset),.clock(clock_27mhz),.noisy(switch[5]),.clean(switch5));
//	debounce sw6(.reset(reset),.clock(clock_27mhz),.noisy(switch[6]),.clean(switch6));
//	debounce sw7(.reset(reset),.clock(clock_27mhz),.noisy(switch[7]),.clean(switch7));
//	debounce bent(.reset(reset),.clock(clock_27mhz),.noisy(~button_enter),.clean(enter));
//   debounce but0(.reset(reset),.clock(clock_27mhz),.noisy(~button0),.clean(b0));
//   debounce but1(.reset(reset),.clock(clock_27mhz),.noisy(~button1),.clean(b1));
//   debounce but2(.reset(reset),.clock(clock_27mhz),.noisy(~button2),.clean(b2));
//   debounce but3(.reset(reset),.clock(clock_27mhz),.noisy(~button3),.clean(b3));
//   debounce butl(.reset(reset),.clock(clock_27mhz),.noisy(~button_left),.clean(bl));
//   debounce butr(.reset(reset),.clock(clock_27mhz),.noisy(~button_right),.clean(br));
//
//	reg [4:0] volume;
//   always @ (posedge clock_27mhz) begin
//     if (reset) volume <= 5'd24;
//     else begin
//	if (vup & ~old_vup & volume != 5'd31) volume <= volume+1;       
//	if (vdown & ~old_vdown & volume != 5'd0) volume <= volume-1;       
//     end
//     old_vup <= vup;
//     old_vdown <= vdown;
//   end
//	wire [17:0] for_ac97_l;
//	wire [17:0] for_ac97_r;
//	wire [9:0] f_controls;
//	wire [9:0] t_controls;
//	wire [10:0] status;
//	wire [55:0] freq_data;
//	
//	// frequency weights output to hex display
//	wire [4:0] test1;
//	wire [4:0] test2;
//	wire [4:0] test3;
//	wire [4:0] test4;
//	wire [4:0] test5;
//	wire [4:0] test6;
//	wire [4:0] test7;
//	
//   //High Level FSM
//	HighLevelFSM HLFSM(.clock(clock_27mhz),.reset(reset),
//							.controls({bl,br,enter,b3,b2,b1,b0,switch7,
//							switch6,switch5,switch4,switch3,switch2,switch1,switch0}),
//							.f_controls(f_controls),.t_controls(t_controls),
//							.status(status));
//	
//	// AC97 driver
//   audio a(clock_27mhz, reset, volume, from_ac97_data_l, for_ac97_l,from_ac97_data_r,for_ac97_r, ready,
//	       audio_reset_b, ac97_sdata_out, ac97_sdata_in,
//	       ac97_synch, ac97_bit_clock);
//	
//	//Assign output data
//	ProcessMod process(.clock(clock_27mhz),.reset(reset),.ready(ready),
//			 .l_audio_in(from_ac97_data_l),.r_audio_in(from_ac97_data_r),
//			 .f_controls(f_controls),.t_controls(t_controls),
//			 .l_audio_out(for_ac97_l),.r_audio_out(for_ac97_r),
//			 .freq1(freq_data[7:0]),.freq2(freq_data[15:8]),
//			 .freq3(freq_data[23:16]),.freq4(freq_data[31:24]),
//			 .freq5(freq_data[39:32]),.freq6(freq_data[47:40]),
//			 .freq7(freq_data[55:48]),.test1(test1),.test2(test2),
//			 .test3(test3),.test4(test4),.test5(test5),.test6(test6),
//			 .test7(test7));
//   
//	display_16hex disp(reset, clock_27mhz,
//			{3'b0,test7,3'b0,test6,3'b0,test5,3'b0,test4,3'b0,test3,
//			3'b0,test2,3'b0,test1}, // bits to output to hex display
//		
//			disp_blank, disp_clock, disp_rs, disp_ce_b,
//			disp_reset_b, disp_data_out);
//	
//	
//	wire [17:0] a_data;
//   wire [29:0] LEDS;
//	assign a_data=for_ac97_l;
//	// show volume during playback.
//   // led is active low
//   assign led = ~{1'b0,status[10],switch0, volume};
//   VDM lights(.clock(clock_27mhz),.reset(reset),.ready(ready),
//              .a_data(a_data[17:0]),.f_data(48'b0),.controls(1'b0),
//              .lights(LEDS));
//
//   assign user4[4:0]=~{LEDS[4:0]};
//   assign user4[12:8]=~{LEDS[9:5]};
//   assign user4[20:16]=~{LEDS[14:10]};
//   assign user3[4:0]=~{LEDS[19:15]};
//   assign user3[12:8]=~{LEDS[24:20]};
//   assign user3[20:16]=~{LEDS[29:25]};
//   // output useful things to the logic analyzer connectors
//   assign analyzer1_clock = ac97_bit_clock;
//   assign analyzer1_data[0] = audio_reset_b;
//   assign analyzer1_data[1] = ac97_sdata_out;
//   assign analyzer1_data[2] = ac97_sdata_in;
//   assign analyzer1_data[3] = ac97_synch;
//   assign analyzer1_data[15:4] = 0;
//
//   assign analyzer3_clock = ready;
//   assign analyzer3_data = {from_ac97_data_l, for_ac97_l};
//endmodule
//
/////////////////////////////////////////////////////////////////////////////////
///// Hex Display Module
/////////////////////////////////////////////////////////////////////////////////
//
//module display_16hex (reset, clock_27mhz, data, 
//		disp_blank, disp_clock, disp_rs, disp_ce_b,
//		disp_reset_b, disp_data_out);
//
//   input reset, clock_27mhz;    // clock and reset (active high reset)
//   input [63:0] data;		// 16 hex nibbles to display
//   
//   output disp_blank, disp_clock, disp_data_out, disp_rs, disp_ce_b, 
//	  disp_reset_b;
//   
//   reg disp_data_out, disp_rs, disp_ce_b, disp_reset_b;
//   
//   ////////////////////////////////////////////////////////////////////////////
//   //
//   // Display Clock
//   //
//   // Generate a 500kHz clock for driving the displays.
//   //
//   ////////////////////////////////////////////////////////////////////////////
//   
//   reg [4:0] count;
//   reg [7:0] reset_count;
//   reg clock;
//   wire dreset;
//
//   always @(posedge clock_27mhz)
//     begin
//	if (reset)
//	  begin
//	     count = 0;
//	     clock = 0;
//	  end
//	else if (count == 26)
//	  begin
//	     clock = ~clock;
//	     count = 5'h00;
//	  end
//	else
//	  count = count+1;
//     end
//   
//   always @(posedge clock_27mhz)
//     if (reset)
//       reset_count <= 100;
//     else
//       reset_count <= (reset_count==0) ? 0 : reset_count-1;
//
//   assign dreset = (reset_count != 0);
//
//   assign disp_clock = ~clock;
//
//   ////////////////////////////////////////////////////////////////////////////
//   //
//   // Display State Machine
//   //
//   ////////////////////////////////////////////////////////////////////////////
//      
//   reg [7:0] state;		// FSM state
//   reg [9:0] dot_index;		// index to current dot being clocked out
//   reg [31:0] control;		// control register
//   reg [3:0] char_index;	// index of current character
//   reg [39:0] dots;		// dots for a single digit 
//   reg [3:0] nibble;		// hex nibble of current character
//   
//   assign disp_blank = 1'b0; // low <= not blanked
//   
//   always @(posedge clock)
//     if (dreset)
//       begin
//	  state <= 0;
//	  dot_index <= 0;
//	  control <= 32'h7F7F7F7F;
//       end
//     else
//       casex (state)
//	 8'h00:
//	   begin
//	      // Reset displays
//	      disp_data_out <= 1'b0; 
//	      disp_rs <= 1'b0; // dot register
//	      disp_ce_b <= 1'b1;
//	      disp_reset_b <= 1'b0;	     
//	      dot_index <= 0;
//	      state <= state+1;
//	   end
//	 
//	 8'h01:
//	   begin
//	      // End reset
//	      disp_reset_b <= 1'b1;
//	      state <= state+1;
//	   end
//	 
//	 8'h02:
//	   begin
//	      // Initialize dot register (set all dots to zero)
//	      disp_ce_b <= 1'b0;
//	      disp_data_out <= 1'b0; // dot_index[0];
//	      if (dot_index == 639)
//		state <= state+1;
//	      else
//		dot_index <= dot_index+1;
//	   end
//	 
//	 8'h03:
//	   begin
//	      // Latch dot data
//	      disp_ce_b <= 1'b1;
//	      dot_index <= 31;		// re-purpose to init ctrl reg
//	      disp_rs <= 1'b1; // Select the control register
//	      state <= state+1;
//	   end
//	 
//	 8'h04:
//	   begin
//	      // Setup the control register
//	      disp_ce_b <= 1'b0;
//	      disp_data_out <= control[31];
//	      control <= {control[30:0], 1'b0};	// shift left
//	      if (dot_index == 0)
//		state <= state+1;
//	      else
//		dot_index <= dot_index-1;
//	   end
//	  
//	 8'h05:
//	   begin
//	      // Latch the control register data / dot data
//	      disp_ce_b <= 1'b1;
//	      dot_index <= 39;		// init for single char
//	      char_index <= 15;		// start with MS char
//	      state <= state+1;
//	      disp_rs <= 1'b0;	 	// Select the dot register
//	   end
//	 
//	 8'h06:
//	   begin
//	      // Load the user's dot data into the dot reg, char by char
//	      disp_ce_b <= 1'b0;
//	      disp_data_out <= dots[dot_index]; // dot data from msb
//	      if (dot_index == 0)
//	        if (char_index == 0)
//	          state <= 5;			// all done, latch data
//		else
//		begin
//		  char_index <= char_index - 1;	// goto next char
//		  dot_index <= 39;
//		end
//	      else
//		dot_index <= dot_index-1;	// else loop thru all dots 
//	   end
//
//       endcase
//
//   always @ (data or char_index)
//     case (char_index)
//       4'h0: 	 	nibble <= data[3:0];
//       4'h1: 	 	nibble <= data[7:4];
//       4'h2: 	 	nibble <= data[11:8];
//       4'h3: 	 	nibble <= data[15:12];
//       4'h4: 	 	nibble <= data[19:16];
//       4'h5: 	 	nibble <= data[23:20];
//       4'h6: 	 	nibble <= data[27:24];
//       4'h7: 	 	nibble <= data[31:28];
//       4'h8: 	 	nibble <= data[35:32];
//       4'h9: 	 	nibble <= data[39:36];
//       4'hA: 	 	nibble <= data[43:40];
//       4'hB: 	 	nibble <= data[47:44];
//       4'hC: 	 	nibble <= data[51:48];
//       4'hD: 	 	nibble <= data[55:52];
//       4'hE: 	 	nibble <= data[59:56];
//       4'hF: 	 	nibble <= data[63:60];
//     endcase
//      
//   always @(nibble)
//     case (nibble)
//       4'h0: dots <= 40'b00111110_01010001_01001001_01000101_00111110;
//       4'h1: dots <= 40'b00000000_01000010_01111111_01000000_00000000;
//       4'h2: dots <= 40'b01100010_01010001_01001001_01001001_01000110;
//       4'h3: dots <= 40'b00100010_01000001_01001001_01001001_00110110;
//       4'h4: dots <= 40'b00011000_00010100_00010010_01111111_00010000;
//       4'h5: dots <= 40'b00100111_01000101_01000101_01000101_00111001;
//       4'h6: dots <= 40'b00111100_01001010_01001001_01001001_00110000;
//       4'h7: dots <= 40'b00000001_01110001_00001001_00000101_00000011;
//       4'h8: dots <= 40'b00110110_01001001_01001001_01001001_00110110;
//       4'h9: dots <= 40'b00000110_01001001_01001001_00101001_00011110;
//       4'hA: dots <= 40'b01111110_00001001_00001001_00001001_01111110;
//       4'hB: dots <= 40'b01111111_01001001_01001001_01001001_00110110;
//       4'hC: dots <= 40'b00111110_01000001_01000001_01000001_00100010;
//       4'hD: dots <= 40'b01111111_01000001_01000001_01000001_00111110;
//       4'hE: dots <= 40'b01111111_01001001_01001001_01001001_01000001;
//       4'hF: dots <= 40'b01111111_00001001_00001001_00001001_00000001;
//     endcase
//   
//endmodule